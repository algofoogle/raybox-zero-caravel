* NGSPICE file created from top_ew_algofoogle.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

.subckt top_ew_algofoogle i_clk i_debug_map_overlay i_debug_trace_overlay i_debug_vec_overlay
+ i_gpout0_sel[0] i_gpout0_sel[1] i_gpout0_sel[2] i_gpout0_sel[3] i_gpout0_sel[4]
+ i_gpout0_sel[5] i_gpout1_sel[0] i_gpout1_sel[1] i_gpout1_sel[2] i_gpout1_sel[3]
+ i_gpout1_sel[4] i_gpout1_sel[5] i_gpout2_sel[0] i_gpout2_sel[1] i_gpout2_sel[2]
+ i_gpout2_sel[3] i_gpout2_sel[4] i_gpout2_sel[5] i_gpout3_sel[0] i_gpout3_sel[1]
+ i_gpout3_sel[2] i_gpout3_sel[3] i_gpout3_sel[4] i_gpout3_sel[5] i_gpout4_sel[0]
+ i_gpout4_sel[1] i_gpout4_sel[2] i_gpout4_sel[3] i_gpout4_sel[4] i_gpout4_sel[5]
+ i_gpout5_sel[0] i_gpout5_sel[1] i_gpout5_sel[2] i_gpout5_sel[3] i_gpout5_sel[4]
+ i_gpout5_sel[5] i_la_invalid i_mode[0] i_mode[1] i_mode[2] i_reg_csb i_reg_mosi
+ i_reg_sclk i_reset_lock_a i_reset_lock_b i_tex_in[0] i_tex_in[1] i_tex_in[2] i_tex_in[3]
+ i_vec_csb i_vec_mosi i_vec_sclk o_gpout[0] o_gpout[1] o_gpout[2] o_gpout[3] o_gpout[4]
+ o_gpout[5] o_hsync o_reset o_rgb[0] o_rgb[10] o_rgb[11] o_rgb[12] o_rgb[13] o_rgb[14]
+ o_rgb[15] o_rgb[16] o_rgb[17] o_rgb[18] o_rgb[19] o_rgb[1] o_rgb[20] o_rgb[21] o_rgb[22]
+ o_rgb[23] o_rgb[2] o_rgb[3] o_rgb[4] o_rgb[5] o_rgb[6] o_rgb[7] o_rgb[8] o_rgb[9]
+ o_tex_csb o_tex_oeb0 o_tex_out0 o_tex_sclk o_vsync ones[0] ones[10] ones[11] ones[12]
+ ones[13] ones[14] ones[15] ones[1] ones[2] ones[3] ones[4] ones[5] ones[6] ones[7]
+ ones[8] ones[9] vccd1 vssd1 zeros[0] zeros[10] zeros[11] zeros[12] zeros[13] zeros[14]
+ zeros[15] zeros[1] zeros[2] zeros[3] zeros[4] zeros[5] zeros[6] zeros[7] zeros[8]
+ zeros[9]
XFILLER_140_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__02438_ clknet_0__02438_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02438_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18869_ _02699_ _03474_ _03462_ _03505_ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__and4b_1
XFILLER_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19025__200 clknet_1_1__leaf__02734_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__inv_2
XFILLER_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19071__242 clknet_1_0__leaf__02738_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__inv_2
XFILLER_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20127_ clknet_leaf_76_i_clk _01058_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09938_ rbzero.tex_r0\[30\] rbzero.tex_r0\[29\] _03017_ vssd1 vssd1 vccd1 vccd1 _03022_
+ sky130_fd_sc_hd__mux2_1
XFILLER_120_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20058_ clknet_leaf_0_i_clk _00989_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.mosi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_09869_ rbzero.tex_r0\[63\] rbzero.tex_r0\[62\] _02984_ vssd1 vssd1 vccd1 vccd1 _02986_
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11900_ _04673_ _04674_ net24 vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__mux2_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12880_ _05634_ _05635_ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__xor2_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ net16 _04603_ _04605_ _04607_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__a31o_1
XFILLER_27_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14550_ _07083_ _07085_ vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__xnor2_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _03782_ _04519_ _04515_ _03865_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__a22o_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13501_ _06103_ _05988_ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__nor2_1
XFILLER_199_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10713_ _03499_ _03500_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__nor2_1
XFILLER_159_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _06759_ _07165_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__or2_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _04473_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__buf_6
X_16220_ _08713_ _08715_ _08711_ vssd1 vssd1 vccd1 vccd1 _08833_ sky130_fd_sc_hd__o21ai_2
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13432_ _06187_ _06182_ _06186_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__and3_1
X_10644_ rbzero.map_overlay.i_otherx\[2\] rbzero.map_rom.f2 vssd1 vssd1 vccd1 vccd1
+ _03440_ sky130_fd_sc_hd__xor2_1
XFILLER_139_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16151_ _08645_ _08655_ _08653_ vssd1 vssd1 vccd1 vccd1 _08764_ sky130_fd_sc_hd__a21o_1
XFILLER_155_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13363_ _06038_ _06065_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__xor2_1
X_10575_ rbzero.debug_overlay.playerX\[3\] _03369_ vssd1 vssd1 vccd1 vccd1 _03371_
+ sky130_fd_sc_hd__or2_1
XFILLER_158_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15102_ _07783_ _07789_ vssd1 vssd1 vccd1 vccd1 _07790_ sky130_fd_sc_hd__nand2_1
XFILLER_6_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12314_ _03480_ _04920_ _05070_ _03489_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__a211oi_2
XFILLER_170_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16082_ _08693_ _08695_ vssd1 vssd1 vccd1 vccd1 _08696_ sky130_fd_sc_hd__xor2_2
X_13294_ _05978_ _06031_ _06049_ _06029_ _06050_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__a221o_1
XFILLER_6_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15033_ _07718_ _07719_ vssd1 vssd1 vccd1 vccd1 _07721_ sky130_fd_sc_hd__and2_1
XFILLER_6_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19910_ clknet_leaf_19_i_clk _00841_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vinf
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_142_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12245_ _04946_ _05006_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__nor2_2
XFILLER_107_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12176_ _03345_ _04923_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__nor2_1
X_19841_ clknet_leaf_15_i_clk _00772_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11127_ _03522_ _03899_ _03912_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__o21ai_4
X_16984_ _09445_ _09450_ _09452_ vssd1 vssd1 vccd1 vccd1 _09590_ sky130_fd_sc_hd__a21oi_1
XFILLER_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19772_ clknet_leaf_6_i_clk _00703_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_95_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18723_ rbzero.debug_overlay.playerY\[-1\] _02582_ _02606_ _02559_ vssd1 vssd1 vccd1
+ vccd1 _01019_ sky130_fd_sc_hd__a211o_1
X_11058_ _03515_ _03344_ _03342_ _03524_ _03843_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__a221o_1
X_15935_ _08524_ _07929_ vssd1 vssd1 vccd1 vccd1 _08554_ sky130_fd_sc_hd__and2_1
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10009_ rbzero.tex_g1\[59\] rbzero.tex_g1\[60\] _02976_ vssd1 vssd1 vccd1 vccd1 _03059_
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18654_ _02534_ _02553_ _02554_ _02356_ vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__o211a_1
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15866_ _08482_ _08481_ _08490_ vssd1 vssd1 vccd1 vccd1 _08494_ sky130_fd_sc_hd__and3_1
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17605_ _01880_ _01884_ _01881_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__a21bo_1
XFILLER_92_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14817_ _06939_ _07157_ vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__nor2_1
XFILLER_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18585_ rbzero.pov.spi_buffer\[60\] rbzero.pov.spi_buffer\[61\] _02510_ vssd1 vssd1
+ vccd1 vccd1 _02512_ sky130_fd_sc_hd__mux2_1
XFILLER_52_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtop_ew_algofoogle_120 vssd1 vssd1 vccd1 vccd1 ones[13] top_ew_algofoogle_120/LO sky130_fd_sc_hd__conb_1
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15797_ rbzero.row_render.texu\[0\] _08456_ _08453_ rbzero.wall_tracer.texu\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__a22o_1
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17536_ rbzero.wall_tracer.rayAddendY\[4\] _01825_ _03509_ vssd1 vssd1 vccd1 vccd1
+ _01826_ sky130_fd_sc_hd__mux2_1
XFILLER_17_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14748_ _06949_ _06966_ _07005_ _07047_ vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__nor4_1
XFILLER_33_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17467_ _01756_ _01760_ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__xnor2_1
X_14679_ _07076_ _07366_ vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__nor2_1
XFILLER_189_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16418_ _09027_ _09028_ vssd1 vssd1 vccd1 vccd1 _09029_ sky130_fd_sc_hd__nand2_1
XFILLER_177_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17398_ rbzero.debug_overlay.playerX\[5\] _01697_ rbzero.wall_tracer.state\[1\] vssd1
+ vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__mux2_1
XFILLER_125_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16349_ rbzero.wall_tracer.trackDistX\[2\] rbzero.wall_tracer.stepDistX\[2\] vssd1
+ vssd1 vccd1 vccd1 _08961_ sky130_fd_sc_hd__or2_1
X_19020__196 clknet_1_0__leaf__02733_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__inv_2
XFILLER_118_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18019_ _02211_ vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09723_ _02901_ _02904_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__and2_1
XFILLER_101_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18389__33 clknet_1_0__leaf__02434_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__inv_2
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10360_ rbzero.tex_b1\[21\] rbzero.tex_b1\[22\] _03243_ vssd1 vssd1 vccd1 vccd1 _03244_
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10291_ _03207_ vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18936__120 clknet_1_1__leaf__02725_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__inv_2
XFILLER_151_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12030_ _04798_ _04799_ _04802_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__a21o_1
XFILLER_105_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13981_ _06727_ vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15720_ _08270_ _08402_ vssd1 vssd1 vccd1 vccd1 _08403_ sky130_fd_sc_hd__xnor2_2
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_52_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_101_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12932_ _05450_ _05688_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__nor2_1
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _07269_ _08333_ vssd1 vssd1 vccd1 vccd1 _08334_ sky130_fd_sc_hd__nor2_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _05433_ _05474_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__or2_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _07262_ _07289_ vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ rbzero.pov.spi_counter\[3\] _02423_ _02425_ _02421_ vssd1 vssd1 vccd1 vccd1
+ _00847_ sky130_fd_sc_hd__o211a_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _03464_ _04566_ _04590_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__a21oi_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _06779_ vssd1 vssd1 vccd1 vccd1 _08266_ sky130_fd_sc_hd__inv_2
XFILLER_187_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12794_ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__clkbuf_4
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_67_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18982__162 clknet_1_0__leaf__02729_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__inv_2
XFILLER_144_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17321_ _01643_ _01644_ _09622_ _01522_ vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__o211a_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _07120_ _07220_ vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__nand2_1
XFILLER_183_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _02981_ _04519_ _04513_ _04521_ _04522_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__a32o_1
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17252_ rbzero.wall_tracer.trackDistY\[-1\] rbzero.wall_tracer.stepDistY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__nor2_1
X_14464_ _04831_ _07149_ _07151_ _03492_ vssd1 vssd1 vccd1 vccd1 _07152_ sky130_fd_sc_hd__a211o_2
X_11676_ _03693_ _04454_ _04456_ _03669_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__o211a_1
XFILLER_186_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16203_ _08786_ _08814_ vssd1 vssd1 vccd1 vccd1 _08816_ sky130_fd_sc_hd__or2_1
X_13415_ _05538_ _06055_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__and2_1
X_19078__248 clknet_1_1__leaf__02739_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__inv_2
X_10627_ rbzero.map_overlay.i_mapdx\[3\] _03413_ _03373_ rbzero.map_overlay.i_mapdx\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__o2bb2a_1
X_17183_ rbzero.wall_tracer.state\[1\] _03493_ _01521_ vssd1 vssd1 vccd1 vccd1 _01526_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_127_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14395_ _07077_ _07079_ _07082_ vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__o21a_1
X_16134_ _07984_ _08081_ vssd1 vssd1 vccd1 vccd1 _08747_ sky130_fd_sc_hd__nor2_1
XFILLER_6_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13346_ _05610_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__clkbuf_4
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10558_ _03353_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__inv_2
XFILLER_183_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16065_ _07199_ _08678_ _08402_ _08400_ vssd1 vssd1 vccd1 vccd1 _08679_ sky130_fd_sc_hd__o31a_1
X_13277_ _06003_ _06033_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__xnor2_4
X_10489_ rbzero.tex_b0\[24\] rbzero.tex_b0\[23\] _03302_ vssd1 vssd1 vccd1 vccd1 _03311_
+ sky130_fd_sc_hd__mux2_1
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15016_ _07272_ _07285_ _07283_ vssd1 vssd1 vccd1 vccd1 _07704_ sky130_fd_sc_hd__a21o_1
XFILLER_130_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12228_ rbzero.wall_tracer.trackDistX\[1\] rbzero.wall_tracer.trackDistY\[1\] vssd1
+ vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__or2b_1
XFILLER_29_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19824_ clknet_leaf_14_i_clk _00755_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12159_ _04886_ _04908_ _04916_ _04920_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__or4b_1
XFILLER_64_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19755_ clknet_leaf_94_i_clk _00686_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16967_ _09570_ _09572_ vssd1 vssd1 vccd1 vccd1 _09573_ sky130_fd_sc_hd__nor2_1
XFILLER_84_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18706_ rbzero.pov.ready_buffer\[47\] _02413_ _02582_ _02594_ vssd1 vssd1 vccd1 vccd1
+ _02595_ sky130_fd_sc_hd__a211o_1
X_15918_ _08524_ _07813_ vssd1 vssd1 vccd1 vccd1 _08539_ sky130_fd_sc_hd__and2_1
X_16898_ _09429_ _09430_ _09504_ vssd1 vssd1 vccd1 vccd1 _09505_ sky130_fd_sc_hd__o21ai_1
X_19686_ clknet_leaf_70_i_clk _00617_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_64_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18637_ _02542_ vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__clkbuf_4
X_15849_ _03369_ _07825_ _08478_ vssd1 vssd1 vccd1 vccd1 _08479_ sky130_fd_sc_hd__a21o_1
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18568_ rbzero.pov.spi_buffer\[52\] rbzero.pov.spi_buffer\[53\] _02499_ vssd1 vssd1
+ vccd1 vccd1 _02503_ sky130_fd_sc_hd__mux2_1
XFILLER_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17519_ _01808_ _01809_ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__nand2_1
X_18499_ rbzero.pov.spi_buffer\[19\] rbzero.pov.spi_buffer\[20\] _02466_ vssd1 vssd1
+ vccd1 vccd1 _02467_ sky130_fd_sc_hd__mux2_1
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20461_ net141 _01392_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19137__301 clknet_1_0__leaf__02745_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__inv_2
XFILLER_146_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20392_ net452 _01323_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19183__343 clknet_1_0__leaf__02749_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__inv_2
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11530_ _03534_ _04309_ _04312_ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__o21a_1
XFILLER_12_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11461_ rbzero.tex_g1\[23\] rbzero.tex_g1\[22\] _03700_ vssd1 vssd1 vccd1 vccd1 _04244_
+ sky130_fd_sc_hd__mux2_1
XFILLER_109_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13200_ _05952_ _05956_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__nor2_1
X_10412_ rbzero.tex_b0\[61\] rbzero.tex_b0\[60\] _03269_ vssd1 vssd1 vccd1 vccd1 _03271_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11392_ rbzero.tex_g0\[15\] rbzero.tex_g0\[14\] _03709_ vssd1 vssd1 vccd1 vccd1 _04176_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14180_ rbzero.wall_tracer.rayAddendY\[-2\] rbzero.wall_tracer.rayAddendX\[-2\] _06849_
+ vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__mux2_1
XFILLER_180_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13131_ _05628_ _05858_ _05887_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__a21o_1
X_10343_ rbzero.tex_b1\[29\] rbzero.tex_b1\[30\] _03232_ vssd1 vssd1 vccd1 vccd1 _03235_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10274_ _03198_ vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__clkbuf_1
X_13062_ _05809_ _05817_ _05818_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__a21oi_1
XFILLER_151_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12013_ _04779_ _04393_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__nor2_1
X_17870_ _02123_ _02127_ _02128_ _02103_ vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__o211a_1
XFILLER_132_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16821_ _09426_ _09427_ vssd1 vssd1 vccd1 vccd1 _09428_ sky130_fd_sc_hd__nor2_1
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16752_ _09133_ _08889_ vssd1 vssd1 vccd1 vccd1 _09360_ sky130_fd_sc_hd__nor2_1
X_19540_ clknet_leaf_38_i_clk _00014_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13964_ rbzero.wall_tracer.stepDistY\[-3\] _06712_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _06713_ sky130_fd_sc_hd__mux2_1
XFILLER_111_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15703_ _08250_ _08378_ _08385_ vssd1 vssd1 vccd1 vccd1 _08386_ sky130_fd_sc_hd__a21o_1
XFILLER_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12915_ _05651_ _05650_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__xnor2_1
X_16683_ _09289_ _09291_ vssd1 vssd1 vccd1 vccd1 _09292_ sky130_fd_sc_hd__xor2_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19471_ clknet_leaf_50_i_clk _00417_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13895_ _06650_ vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15634_ _08316_ vssd1 vssd1 vccd1 vccd1 _08317_ sky130_fd_sc_hd__clkbuf_4
XFILLER_46_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12846_ _05600_ _05601_ _05602_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__o21ba_1
XFILLER_34_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _02412_ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__clkbuf_4
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _06970_ _07748_ vssd1 vssd1 vccd1 vccd1 _08249_ sky130_fd_sc_hd__or2_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _05210_ _05424_ _05417_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__and3_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _01622_ _01624_ _01623_ vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__o21ba_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _07192_ _07202_ vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__nor2_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11728_ net4 _04502_ _04505_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__nand3_1
X_18284_ _02374_ vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__clkbuf_1
X_15496_ _07827_ _08179_ _04832_ vssd1 vssd1 vccd1 vccd1 _08181_ sky130_fd_sc_hd__a21o_1
XFILLER_174_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17235_ _01569_ _01570_ _01558_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__o21ai_1
X_14447_ _06860_ rbzero.wall_tracer.stepDistY\[1\] _04840_ vssd1 vssd1 vccd1 vccd1
+ _07135_ sky130_fd_sc_hd__o21ai_1
X_11659_ _03656_ _04437_ _04438_ _04439_ _03673_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__o221a_1
XFILLER_174_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17166_ _01474_ _01509_ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__xnor2_2
X_14378_ _06865_ _07052_ vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__or2_1
XFILLER_183_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16117_ _07856_ _08191_ vssd1 vssd1 vccd1 vccd1 _08730_ sky130_fd_sc_hd__nor2_1
X_13329_ _05768_ _06055_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__and2_1
X_17097_ _09700_ _09701_ vssd1 vssd1 vccd1 vccd1 _09702_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1__f__02755_ clknet_0__02755_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02755_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16048_ _08265_ _08392_ _08393_ _08389_ vssd1 vssd1 vccd1 vccd1 _08662_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19807_ clknet_leaf_2_i_clk _00738_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17999_ rbzero.pov.spi_buffer\[52\] rbzero.pov.ready_buffer\[52\] _02197_ vssd1 vssd1
+ vccd1 vccd1 _02201_ sky130_fd_sc_hd__mux2_1
XFILLER_78_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18989__168 clknet_1_1__leaf__02730_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__inv_2
X_19738_ clknet_leaf_91_i_clk _00669_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19669_ clknet_leaf_11_i_clk _00600_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f2 sky130_fd_sc_hd__dfxtp_1
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18906__93 clknet_1_1__leaf__02441_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__inv_2
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20513_ clknet_leaf_78_i_clk _01444_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20444_ net504 _01375_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20375_ net435 _01306_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10961_ rbzero.tex_r0\[57\] rbzero.tex_r0\[56\] _03663_ vssd1 vssd1 vccd1 vccd1 _03747_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12700_ _05356_ _05456_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__nand2_1
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13680_ _06421_ _06420_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__and2b_1
X_10892_ _03675_ _03676_ _03677_ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__mux2_1
XFILLER_43_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12631_ _05385_ _05387_ _05380_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__mux2_1
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15350_ _07991_ _08035_ vssd1 vssd1 vccd1 vccd1 _08036_ sky130_fd_sc_hd__xnor2_2
XFILLER_12_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12562_ _05318_ _05246_ _05251_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__and3b_1
XFILLER_15_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14301_ _06987_ _06988_ vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__nand2_1
X_11513_ _04293_ _04294_ _04295_ _03726_ _03689_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__o221a_1
X_15281_ _07790_ _07844_ vssd1 vssd1 vccd1 vccd1 _07967_ sky130_fd_sc_hd__nor2_1
XFILLER_184_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12493_ _05221_ _05222_ _05223_ _05249_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__or4_1
X_17020_ _09623_ _09624_ _09625_ vssd1 vssd1 vccd1 vccd1 _09626_ sky130_fd_sc_hd__a21oi_1
X_14232_ _06919_ _06899_ _06917_ vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__or3_2
XFILLER_172_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11444_ _04225_ _04227_ net41 _03541_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__o211a_1
XFILLER_184_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14163_ _06851_ _03496_ _06788_ _03498_ vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__o211a_1
X_11375_ _03740_ _04154_ _04157_ _04158_ _03702_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__o221a_1
XFILLER_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13114_ _05864_ _05869_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__nand2_1
X_10326_ rbzero.tex_b1\[37\] rbzero.tex_b1\[38\] _03221_ vssd1 vssd1 vccd1 vccd1 _03226_
+ sky130_fd_sc_hd__mux2_1
XFILLER_98_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14094_ rbzero.wall_tracer.trackDistY\[7\] _06785_ _06810_ vssd1 vssd1 vccd1 vccd1
+ _00446_ sky130_fd_sc_hd__o21a_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17922_ _02160_ vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__clkbuf_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _05774_ _05787_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__xor2_1
XFILLER_112_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10257_ rbzero.tex_g0\[7\] rbzero.tex_g0\[6\] _03188_ vssd1 vssd1 vccd1 vccd1 _03190_
+ sky130_fd_sc_hd__mux2_1
XFILLER_105_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10188_ _03153_ vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__clkbuf_1
X_17853_ rbzero.spi_registers.spi_counter\[3\] _01660_ _02111_ _02113_ vssd1 vssd1
+ vccd1 vccd1 _02114_ sky130_fd_sc_hd__nor4_1
XFILLER_182_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16804_ _09305_ _09303_ _09302_ vssd1 vssd1 vccd1 vccd1 _09412_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14996_ _07665_ _07682_ _07683_ _07676_ _07681_ vssd1 vssd1 vccd1 vccd1 _07684_ sky130_fd_sc_hd__o32a_1
X_17784_ _02000_ rbzero.wall_tracer.rayAddendX\[6\] vssd1 vssd1 vccd1 vccd1 _02050_
+ sky130_fd_sc_hd__xor2_1
XFILLER_81_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19523_ clknet_leaf_49_i_clk _00469_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[8\]
+ sky130_fd_sc_hd__dfxtp_2
X_16735_ _09341_ _09336_ vssd1 vssd1 vccd1 vccd1 _09343_ sky130_fd_sc_hd__and2b_1
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13947_ _05325_ _06635_ _05271_ vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__a21o_1
XFILLER_19_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16666_ _09273_ _09274_ vssd1 vssd1 vccd1 vccd1 _09275_ sky130_fd_sc_hd__and2_1
X_19454_ clknet_leaf_69_i_clk _00012_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rcp_sel\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_13878_ _05324_ _06595_ _06597_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__and3_1
XFILLER_90_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15617_ _08064_ _08062_ vssd1 vssd1 vccd1 vccd1 _08301_ sky130_fd_sc_hd__nand2_1
XFILLER_22_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12829_ _05583_ _05585_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__xnor2_1
X_16597_ _09107_ _09108_ vssd1 vssd1 vccd1 vccd1 _09206_ sky130_fd_sc_hd__or2b_1
X_19385_ _02859_ _02860_ _02861_ _02854_ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__a22o_1
XFILLER_201_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15548_ _08230_ _08231_ vssd1 vssd1 vccd1 vccd1 _08232_ sky130_fd_sc_hd__nand2_1
X_18336_ _02403_ vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__clkbuf_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18267_ rbzero.spi_registers.spi_buffer\[3\] rbzero.spi_registers.new_sky\[3\] _02361_
+ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__mux2_1
X_15479_ _07991_ _08035_ _08163_ vssd1 vssd1 vccd1 vccd1 _08164_ sky130_fd_sc_hd__a21oi_2
XFILLER_30_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17218_ _01553_ _01554_ _01555_ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__a21oi_1
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18198_ rbzero.spi_registers.new_leak\[5\] _02310_ _02318_ _02314_ vssd1 vssd1 vccd1
+ vccd1 _00782_ sky130_fd_sc_hd__o211a_1
XFILLER_129_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17149_ _01488_ _01492_ vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20160_ net220 _01091_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[7\] sky130_fd_sc_hd__dfxtp_1
X_09971_ _02983_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__clkbuf_4
XFILLER_170_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__02738_ clknet_0__02738_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02738_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20091_ clknet_leaf_8_i_clk _01022_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_85_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20427_ net487 _01358_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11160_ rbzero.tex_r1\[43\] _03664_ _03944_ _03677_ vssd1 vssd1 vccd1 vccd1 _03945_
+ sky130_fd_sc_hd__o211a_1
X_20358_ net418 _01289_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10111_ rbzero.tex_g1\[11\] rbzero.tex_g1\[12\] _03106_ vssd1 vssd1 vccd1 vccd1 _03113_
+ sky130_fd_sc_hd__mux2_1
X_11091_ rbzero.map_overlay.i_otherx\[1\] _03463_ _03466_ _03872_ _03876_ vssd1 vssd1
+ vccd1 vccd1 _03877_ sky130_fd_sc_hd__a221o_1
X_20289_ net349 _01220_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10042_ rbzero.tex_g1\[44\] rbzero.tex_g1\[45\] _03073_ vssd1 vssd1 vccd1 vccd1 _03077_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14850_ _07489_ _07537_ vssd1 vssd1 vccd1 vccd1 _07538_ sky130_fd_sc_hd__xor2_1
XFILLER_75_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13801_ _06474_ _06509_ _06510_ _06557_ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__a22o_1
XFILLER_152_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14781_ _07444_ _07467_ vssd1 vssd1 vccd1 vccd1 _07469_ sky130_fd_sc_hd__nor2_1
XFILLER_112_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11993_ net30 _04742_ _04763_ _04764_ _04766_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__a311o_1
XFILLER_57_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16520_ _09098_ _09129_ vssd1 vssd1 vccd1 vccd1 _09130_ sky130_fd_sc_hd__xnor2_1
XFILLER_28_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13732_ _05551_ _06155_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__or2_1
X_10944_ _03697_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__buf_4
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18440__79 clknet_1_0__leaf__02439_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__inv_2
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16451_ _08908_ _08937_ _08935_ vssd1 vssd1 vccd1 vccd1 _09062_ sky130_fd_sc_hd__a21oi_1
X_13663_ _06400_ _06401_ _06419_ vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__a21o_1
X_10875_ _03660_ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__buf_4
XFILLER_32_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15402_ _08075_ _08086_ vssd1 vssd1 vccd1 vccd1 _08087_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12614_ _05116_ _05311_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__nand2_1
X_16382_ _08991_ _08992_ vssd1 vssd1 vccd1 vccd1 _08993_ sky130_fd_sc_hd__and2b_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13594_ _06343_ _06350_ vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__or2_1
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18121_ rbzero.spi_registers.new_other\[9\] _02264_ _02270_ _02266_ vssd1 vssd1 vccd1
+ vccd1 _00753_ sky130_fd_sc_hd__o211a_1
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15333_ _07199_ _08018_ vssd1 vssd1 vccd1 vccd1 _08019_ sky130_fd_sc_hd__nor2_1
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12545_ _05234_ _05238_ _05275_ _05246_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__o31ai_4
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18052_ rbzero.spi_registers.spi_buffer\[2\] rbzero.spi_registers.spi_buffer\[1\]
+ _02227_ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__mux2_1
X_15264_ _07837_ _07840_ _07836_ vssd1 vssd1 vccd1 vccd1 _07950_ sky130_fd_sc_hd__a21bo_1
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12476_ _05220_ _05224_ _05226_ _05232_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__or4_1
X_17003_ _09426_ _09608_ vssd1 vssd1 vccd1 vccd1 _09609_ sky130_fd_sc_hd__nand2_1
XFILLER_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14215_ _04907_ _05091_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__mux2_1
X_11427_ rbzero.tex_g0\[39\] rbzero.tex_g0\[38\] _03614_ vssd1 vssd1 vccd1 vccd1 _04211_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_5 _04307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15195_ _07733_ _07880_ _07881_ vssd1 vssd1 vccd1 vccd1 _07882_ sky130_fd_sc_hd__o21ai_1
XFILLER_99_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14146_ rbzero.wall_tracer.stepDistX\[10\] _06781_ _04833_ vssd1 vssd1 vccd1 vccd1
+ _06838_ sky130_fd_sc_hd__mux2_1
X_11358_ rbzero.debug_overlay.playerY\[-1\] _04093_ _04137_ _04142_ vssd1 vssd1 vccd1
+ vccd1 _04143_ sky130_fd_sc_hd__a211o_1
XFILLER_99_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10309_ rbzero.tex_b1\[45\] rbzero.tex_b1\[46\] _03210_ vssd1 vssd1 vccd1 vccd1 _03217_
+ sky130_fd_sc_hd__mux2_1
XFILLER_193_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18954_ clknet_1_1__leaf__02440_ vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__buf_1
X_14077_ rbzero.wall_tracer.visualWallDist\[-1\] _06796_ _06791_ rbzero.wall_tracer.trackDistX\[-1\]
+ _06797_ vssd1 vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__o221a_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11289_ _04046_ _04057_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__or2_1
XFILLER_140_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17905_ _02151_ vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__clkbuf_1
X_13028_ _05784_ _05782_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18885_ _04508_ _02709_ _02711_ _02285_ vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__a22o_1
XFILLER_121_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17836_ _02001_ rbzero.wall_tracer.rayAddendX\[10\] vssd1 vssd1 vccd1 vccd1 _02098_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17767_ _02030_ _02031_ _03339_ _02034_ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_35_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14979_ _07650_ _07666_ vssd1 vssd1 vccd1 vccd1 _07667_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19506_ clknet_leaf_55_i_clk _00452_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
X_16718_ _08000_ _07993_ _07960_ _08070_ vssd1 vssd1 vccd1 vccd1 _09326_ sky130_fd_sc_hd__or4_1
X_17698_ _08458_ _01965_ _01966_ _01970_ vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__a31o_1
XFILLER_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19437_ _02889_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16649_ _09255_ _09257_ vssd1 vssd1 vccd1 vccd1 _09258_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19368_ _02846_ _02847_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18319_ rbzero.spi_registers.new_other\[6\] rbzero.spi_registers.spi_buffer\[6\]
+ _02388_ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__mux2_1
XFILLER_187_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19299_ _02785_ _02786_ _02788_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__o21ai_1
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20212_ net272 _01143_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20143_ clknet_leaf_12_i_clk _01074_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[1\] sky130_fd_sc_hd__dfxtp_2
X_09954_ _03030_ vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20074_ clknet_leaf_86_i_clk _01005_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_09885_ rbzero.tex_r0\[55\] rbzero.tex_r0\[54\] _02984_ vssd1 vssd1 vccd1 vccd1 _02994_
+ sky130_fd_sc_hd__mux2_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18930__115 clknet_1_1__leaf__02724_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__inv_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10660_ _03409_ _03419_ _03429_ _03455_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__or4b_1
XFILLER_179_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10591_ rbzero.wall_tracer.visualWallDist\[9\] rbzero.wall_tracer.visualWallDist\[8\]
+ _03384_ _03386_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__or4_1
XFILLER_167_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12330_ _03488_ _05086_ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__nand2_1
XFILLER_182_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12261_ rbzero.wall_tracer.mapY\[9\] _04929_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__xnor2_1
XFILLER_182_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14000_ _06603_ _06634_ _06728_ _05315_ vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__a22o_1
X_11212_ rbzero.row_render.side _03631_ rbzero.row_render.wall\[0\] vssd1 vssd1 vccd1
+ vccd1 _03997_ sky130_fd_sc_hd__a21oi_1
XFILLER_107_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12192_ rbzero.wall_tracer.trackDistY\[9\] vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__inv_2
XFILLER_134_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11143_ rbzero.tex_r1\[48\] _03920_ _03925_ _03927_ vssd1 vssd1 vccd1 vccd1 _03928_
+ sky130_fd_sc_hd__a31o_1
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 o_rgb[22] sky130_fd_sc_hd__buf_2
XFILLER_122_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11074_ _03851_ _03853_ _03859_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__and3_1
X_15951_ rbzero.wall_tracer.trackDistX\[-4\] _08553_ _08561_ _08568_ vssd1 vssd1 vccd1
+ vccd1 _00545_ sky130_fd_sc_hd__o22a_1
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10025_ _03067_ vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__clkbuf_1
X_14902_ _06969_ _06977_ _07157_ _07178_ vssd1 vssd1 vccd1 vccd1 _07590_ sky130_fd_sc_hd__or4_1
X_18670_ rbzero.debug_overlay.playerX\[2\] rbzero.debug_overlay.playerX\[1\] _02561_
+ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__or3_1
X_15882_ _08506_ vssd1 vssd1 vccd1 vccd1 _08507_ sky130_fd_sc_hd__buf_4
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17621_ _01901_ _03345_ _05009_ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__mux2_1
X_14833_ _07517_ _07519_ _07520_ vssd1 vssd1 vccd1 vccd1 _07521_ sky130_fd_sc_hd__a21oi_1
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ rbzero.wall_tracer.rayAddendY\[5\] _08447_ _01840_ _01714_ vssd1 vssd1 vccd1
+ vccd1 _01841_ sky130_fd_sc_hd__a22o_1
X_14764_ _06908_ _07177_ _07450_ _07451_ _07384_ vssd1 vssd1 vccd1 vccd1 _07452_ sky130_fd_sc_hd__o32a_1
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ net27 vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__buf_2
XFILLER_189_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16503_ _07878_ _07787_ _08987_ vssd1 vssd1 vccd1 vccd1 _09113_ sky130_fd_sc_hd__or3_1
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13715_ _06430_ _06471_ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__xnor2_1
X_10927_ _03710_ _03711_ _03712_ _03666_ _03670_ vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__o221a_1
XFILLER_32_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17483_ _01759_ _01774_ _01773_ _01772_ vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__o211ai_2
XFILLER_45_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14695_ _07345_ _07382_ vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__xnor2_1
XFILLER_189_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16434_ _09031_ _09044_ vssd1 vssd1 vccd1 vccd1 _09045_ sky130_fd_sc_hd__xor2_2
X_13646_ _06373_ _06363_ _06372_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__nand3_1
X_10858_ _03638_ _03641_ rbzero.row_render.side vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__o21ai_1
XFILLER_176_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _08107_ _07984_ _07960_ _08070_ vssd1 vssd1 vccd1 vccd1 _08976_ sky130_fd_sc_hd__or4_1
XFILLER_158_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13577_ _06286_ _06329_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__and2_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10789_ rbzero.texV\[8\] _03573_ _03574_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__a21boi_1
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15316_ _07999_ _08001_ vssd1 vssd1 vccd1 vccd1 _08002_ sky130_fd_sc_hd__xnor2_1
X_18104_ _03906_ vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__inv_2
XFILLER_185_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12528_ _05235_ _05276_ _05284_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__and3_1
X_16296_ _08883_ _08907_ vssd1 vssd1 vccd1 vccd1 _08908_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18035_ _02219_ vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__clkbuf_1
X_15247_ _07810_ _07822_ _07933_ vssd1 vssd1 vccd1 vccd1 _07934_ sky130_fd_sc_hd__a21o_1
XFILLER_173_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12459_ _05199_ _05127_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__nand2_1
XFILLER_132_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15178_ _07235_ vssd1 vssd1 vccd1 vccd1 _07865_ sky130_fd_sc_hd__clkbuf_4
XFILLER_99_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14129_ _06829_ vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19986_ clknet_leaf_95_i_clk _00917_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__02437_ clknet_0__02437_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02437_
+ sky130_fd_sc_hd__clkbuf_16
X_18868_ _03865_ _03459_ _02903_ _03529_ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__or4_1
XFILLER_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17819_ _02001_ _01972_ _02082_ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__a21oi_1
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18799_ rbzero.pov.ready_buffer\[27\] _02636_ _02659_ _02643_ vssd1 vssd1 vccd1 vccd1
+ _01042_ sky130_fd_sc_hd__o211a_1
XFILLER_36_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09937_ _03021_ vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20126_ clknet_leaf_91_i_clk _01057_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20057_ clknet_leaf_7_i_clk _00988_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[73\]
+ sky130_fd_sc_hd__dfxtp_1
X_09868_ _02985_ vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__clkbuf_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _02947_ vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__clkbuf_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ net16 _04606_ _04584_ net20 net19 vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__o2111ai_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _04522_ _04528_ _04531_ _04538_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__a211o_1
XFILLER_198_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13500_ _06168_ _06256_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__xnor2_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__inv_2
XFILLER_187_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _07157_ _07158_ _07167_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__nor3_2
XFILLER_187_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _04471_ _04472_ _04148_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__o21a_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ _06182_ _06186_ _06187_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__a21oi_1
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10643_ rbzero.map_overlay.i_otherx\[4\] _03364_ _03390_ _03437_ _03438_ vssd1 vssd1
+ vccd1 vccd1 _03439_ sky130_fd_sc_hd__a221o_1
XFILLER_139_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16150_ _08728_ _08762_ vssd1 vssd1 vccd1 vccd1 _08763_ sky130_fd_sc_hd__xnor2_1
XFILLER_167_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13362_ _06100_ _06101_ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10574_ rbzero.debug_overlay.playerX\[3\] _03369_ vssd1 vssd1 vccd1 vccd1 _03370_
+ sky130_fd_sc_hd__nand2_1
XFILLER_155_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15101_ _07785_ _07788_ vssd1 vssd1 vccd1 vccd1 _07789_ sky130_fd_sc_hd__nor2_1
XFILLER_166_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12313_ rbzero.wall_tracer.visualWallDist\[1\] _03480_ vssd1 vssd1 vccd1 vccd1 _05070_
+ sky130_fd_sc_hd__nor2_1
XFILLER_182_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16081_ _08388_ _08410_ _08694_ vssd1 vssd1 vccd1 vccd1 _08695_ sky130_fd_sc_hd__a21oi_2
XFILLER_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13293_ _06029_ _06049_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__nor2_1
XFILLER_6_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15032_ _07718_ _07719_ vssd1 vssd1 vccd1 vccd1 _07720_ sky130_fd_sc_hd__nor2_1
X_12244_ _04951_ _04952_ _05005_ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__or3b_4
XFILLER_107_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19840_ clknet_leaf_15_i_clk _00771_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12175_ _03346_ _04928_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__nor2_1
XFILLER_69_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11126_ _03522_ _03905_ _03910_ _03911_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__a211oi_4
X_19771_ clknet_leaf_6_i_clk _00702_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_16983_ _09578_ _09588_ vssd1 vssd1 vccd1 vccd1 _09589_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18722_ rbzero.pov.ready_buffer\[52\] _02411_ _02535_ _07028_ _02587_ vssd1 vssd1
+ vccd1 vccd1 _02606_ sky130_fd_sc_hd__o221a_1
X_11057_ rbzero.debug_overlay.playerX\[1\] _03463_ _03838_ _03839_ _03842_ vssd1 vssd1
+ vccd1 vccd1 _03843_ sky130_fd_sc_hd__a221o_1
X_15934_ _08507_ vssd1 vssd1 vccd1 vccd1 _08553_ sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10008_ _03058_ vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18653_ _06990_ _02533_ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__nand2_1
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15865_ rbzero.wall_tracer.mapX\[8\] _07826_ vssd1 vssd1 vccd1 vccd1 _08493_ sky130_fd_sc_hd__xor2_1
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17604_ _01757_ _01875_ _03339_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__o21ai_1
XFILLER_149_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14816_ _06969_ _07148_ vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__nor2_1
X_18584_ _02511_ vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__clkbuf_1
Xtop_ew_algofoogle_110 vssd1 vssd1 vccd1 vccd1 ones[3] top_ew_algofoogle_110/LO sky130_fd_sc_hd__conb_1
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15796_ rbzero.row_render.size\[10\] _08456_ _06746_ _08455_ vssd1 vssd1 vccd1 vccd1
+ _00502_ sky130_fd_sc_hd__a22o_1
Xtop_ew_algofoogle_121 vssd1 vssd1 vccd1 vccd1 ones[14] top_ew_algofoogle_121/LO sky130_fd_sc_hd__conb_1
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17535_ _01816_ _01817_ _01824_ _03484_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__o22a_1
X_11959_ _03464_ _04724_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__and2_1
X_14747_ _06966_ _07047_ vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__or2_1
XFILLER_178_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14678_ _06876_ _07075_ vssd1 vssd1 vccd1 vccd1 _07366_ sky130_fd_sc_hd__and2_1
XFILLER_33_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17466_ _01758_ _01759_ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__or2_1
XFILLER_177_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16417_ _08917_ _08920_ _09026_ vssd1 vssd1 vccd1 vccd1 _09028_ sky130_fd_sc_hd__nand3_1
X_13629_ _05697_ _06055_ _06384_ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__a21o_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17397_ _08468_ _01696_ vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16348_ rbzero.wall_tracer.trackDistX\[2\] rbzero.wall_tracer.stepDistX\[2\] vssd1
+ vssd1 vccd1 vccd1 _08960_ sky130_fd_sc_hd__nand2_1
XFILLER_185_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16279_ _08887_ _08890_ vssd1 vssd1 vccd1 vccd1 _08891_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19055__227 clknet_1_1__leaf__02737_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__inv_2
X_18018_ rbzero.pov.spi_buffer\[61\] rbzero.pov.ready_buffer\[61\] _02208_ vssd1 vssd1
+ vccd1 vccd1 _02211_ sky130_fd_sc_hd__mux2_1
XFILLER_145_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19969_ net198 _00900_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09722_ _02902_ _02903_ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__nor2_1
XFILLER_86_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10290_ rbzero.tex_b1\[54\] rbzero.tex_b1\[55\] _03199_ vssd1 vssd1 vccd1 vccd1 _03207_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20109_ clknet_leaf_76_i_clk _01040_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-6\]
+ sky130_fd_sc_hd__dfxtp_2
X_13980_ rbzero.wall_tracer.stepDistY\[-1\] _06726_ _06718_ vssd1 vssd1 vccd1 vccd1
+ _06727_ sky130_fd_sc_hd__mux2_1
XFILLER_58_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12931_ _05655_ _05657_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__xnor2_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15650_ _08191_ vssd1 vssd1 vccd1 vccd1 _08333_ sky130_fd_sc_hd__clkbuf_4
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ _05618_ _05606_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__nand2_1
XFILLER_74_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _07287_ _07288_ vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__nand2_1
XFILLER_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11813_ _03474_ _04569_ _04589_ net17 vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__a211o_1
XFILLER_160_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15581_ _07673_ _08144_ vssd1 vssd1 vccd1 vccd1 _08265_ sky130_fd_sc_hd__nand2_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19160__322 clknet_1_0__leaf__02747_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__inv_2
X_12793_ _05488_ _05489_ _05490_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__nor3_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14532_ _06893_ _07092_ vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__or2_1
X_17320_ _01640_ _01641_ _01642_ _03341_ vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__a31o_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ net6 net5 vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__and2b_1
XFILLER_144_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _06850_ _04886_ _07150_ _06853_ vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__o211a_1
X_17251_ _04964_ _07115_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__nor2_1
XFILLER_109_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11675_ _03823_ _04455_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__or2_1
XFILLER_30_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16202_ _08786_ _08814_ vssd1 vssd1 vccd1 vccd1 _08815_ sky130_fd_sc_hd__nand2_1
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13414_ _06123_ _06128_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__xor2_1
X_10626_ _03420_ _03421_ rbzero.map_rom.i_col\[4\] vssd1 vssd1 vccd1 vccd1 _03422_
+ sky130_fd_sc_hd__a21o_1
X_17182_ rbzero.wall_tracer.trackDistY\[-11\] rbzero.wall_tracer.stepDistY\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__or2_1
XFILLER_168_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14394_ _07080_ _07081_ vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__nand2_1
X_16133_ _08743_ _08744_ _08745_ vssd1 vssd1 vccd1 vccd1 _08746_ sky130_fd_sc_hd__o21a_1
X_13345_ _06100_ _06101_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__nand2_1
X_10557_ rbzero.map_rom.f2 vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__clkbuf_4
XFILLER_6_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16064_ _04841_ rbzero.wall_tracer.stepDistX\[9\] _08269_ _08677_ vssd1 vssd1 vccd1
+ vccd1 _08678_ sky130_fd_sc_hd__a2bb2o_4
X_13276_ _06004_ _06032_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__xnor2_4
XFILLER_182_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10488_ _03310_ vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15015_ _07372_ _07478_ _07700_ _07702_ vssd1 vssd1 vccd1 vccd1 _07703_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_190_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12227_ rbzero.wall_tracer.trackDistX\[-3\] _04986_ _04970_ rbzero.wall_tracer.trackDistX\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__o22a_1
XFILLER_155_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19823_ clknet_leaf_14_i_clk _00754_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12158_ _04917_ _04919_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__xnor2_1
XFILLER_150_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11109_ _03847_ _03894_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__nor2_1
XFILLER_111_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19754_ clknet_leaf_88_i_clk _00685_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16966_ _07993_ _08333_ _09434_ _09571_ vssd1 vssd1 vccd1 vccd1 _09572_ sky130_fd_sc_hd__o31a_1
X_12089_ rbzero.debug_overlay.facingY\[-5\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__nor2_1
XFILLER_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18705_ _06924_ _02535_ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__nor2_1
X_15917_ rbzero.wall_tracer.trackDistX\[-8\] _08508_ _08532_ _08538_ vssd1 vssd1 vccd1
+ vccd1 _00541_ sky130_fd_sc_hd__o22a_1
X_19685_ clknet_leaf_68_i_clk _00616_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16897_ _09464_ _09503_ vssd1 vssd1 vccd1 vccd1 _09504_ sky130_fd_sc_hd__xnor2_1
X_18636_ net39 _02532_ _02261_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__o21a_2
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15848_ _08474_ _08477_ _08475_ vssd1 vssd1 vccd1 vccd1 _08478_ sky130_fd_sc_hd__a21bo_1
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18567_ _02502_ vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15779_ rbzero.wall_tracer.state\[14\] _03484_ _08450_ vssd1 vssd1 vccd1 vccd1 _08451_
+ sky130_fd_sc_hd__and3_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11708__1 clknet_1_1__leaf__04486_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__inv_2
X_17518_ _04109_ rbzero.debug_overlay.vplaneY\[-6\] _01807_ vssd1 vssd1 vccd1 vccd1
+ _01809_ sky130_fd_sc_hd__o21ai_1
XFILLER_33_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18498_ _02443_ vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__clkbuf_4
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17449_ rbzero.wall_tracer.rayAddendY\[-2\] _00013_ _01741_ _01744_ vssd1 vssd1 vccd1
+ vccd1 _00607_ sky130_fd_sc_hd__o22a_1
XFILLER_162_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20460_ net140 _01391_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[51\] sky130_fd_sc_hd__dfxtp_1
X_20391_ net451 _01322_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18966__147 clknet_1_0__leaf__02728_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__inv_2
XFILLER_83_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11460_ rbzero.tex_g1\[21\] rbzero.tex_g1\[20\] _03700_ vssd1 vssd1 vccd1 vccd1 _04243_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19003__181 clknet_1_1__leaf__02731_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__inv_2
X_10411_ _03270_ vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11391_ _04171_ _04174_ _03702_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__mux2_1
XFILLER_136_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13130_ _05875_ _05886_ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__xnor2_1
X_10342_ _03234_ vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13061_ _05783_ _05785_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__xnor2_1
X_10273_ rbzero.tex_b1\[62\] rbzero.tex_b1\[63\] _03117_ vssd1 vssd1 vccd1 vccd1 _03198_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19247__21 clknet_1_0__leaf__02755_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__inv_2
X_12012_ net37 _04783_ _04784_ net36 vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__a31o_1
XFILLER_78_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16820_ _09351_ _09424_ _09425_ vssd1 vssd1 vccd1 vccd1 _09427_ sky130_fd_sc_hd__and3_1
XFILLER_78_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16751_ _09357_ _09358_ vssd1 vssd1 vccd1 vccd1 _09359_ sky130_fd_sc_hd__nand2_1
XFILLER_19_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13963_ _06707_ _06637_ _06711_ _05476_ _06629_ vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__a221o_2
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15702_ _08379_ _08384_ vssd1 vssd1 vccd1 vccd1 _08385_ sky130_fd_sc_hd__xnor2_1
X_12914_ _05666_ _05670_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__xor2_1
X_19470_ clknet_leaf_52_i_clk _00416_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16682_ _09153_ _09174_ _09290_ vssd1 vssd1 vccd1 vccd1 _09291_ sky130_fd_sc_hd__a21oi_2
XFILLER_59_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13894_ rbzero.wall_tracer.stepDistY\[-10\] _06649_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _06650_ sky130_fd_sc_hd__mux2_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15633_ rbzero.wall_tracer.visualWallDist\[10\] _07256_ vssd1 vssd1 vccd1 vccd1 _08316_
+ sky130_fd_sc_hd__and2_1
X_12845_ _05599_ _05574_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__and2b_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _02261_ _02411_ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__nand2_2
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _08247_ _08130_ vssd1 vssd1 vccd1 vccd1 _08248_ sky130_fd_sc_hd__nor2_1
XFILLER_15_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12776_ _05524_ _05532_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__or2_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ rbzero.wall_tracer.trackDistY\[6\] rbzero.wall_tracer.stepDistY\[6\] vssd1
+ vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__and2_1
XFILLER_42_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11727_ _03852_ _04487_ _04496_ _04504_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__a211o_1
X_14515_ _07192_ _07202_ vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__xor2_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ _07827_ _08179_ vssd1 vssd1 vccd1 vccd1 _08180_ sky130_fd_sc_hd__nor2_1
X_18283_ rbzero.spi_registers.spi_buffer\[3\] rbzero.spi_registers.new_floor\[3\]
+ _02370_ vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__mux2_1
XFILLER_187_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17234_ _01566_ _01567_ _01568_ _04946_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__a31o_1
X_11658_ rbzero.tex_b1\[26\] _03690_ _03823_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__a21o_1
X_14446_ _04831_ _07131_ _07133_ vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__a21oi_2
XFILLER_128_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10609_ _03395_ _03390_ _03399_ _03403_ _03404_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__o311a_1
X_17165_ _01476_ _01508_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__xnor2_1
X_14377_ _07055_ _07058_ vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11589_ rbzero.tex_b0\[15\] _04155_ _04156_ _03611_ vssd1 vssd1 vccd1 vccd1 _04371_
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16116_ _08659_ _08637_ vssd1 vssd1 vccd1 vccd1 _08729_ sky130_fd_sc_hd__or2b_1
XFILLER_143_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13328_ _06080_ _06081_ _06084_ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__a21o_1
XFILLER_171_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17096_ _09630_ _09604_ _09699_ vssd1 vssd1 vccd1 vccd1 _09701_ sky130_fd_sc_hd__and3_1
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__02754_ clknet_0__02754_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02754_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16047_ _08249_ _08382_ _08381_ vssd1 vssd1 vccd1 vccd1 _08661_ sky130_fd_sc_hd__o21ba_1
X_13259_ _06015_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__inv_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19806_ clknet_leaf_2_i_clk _00737_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_97_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17998_ _02200_ vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__clkbuf_1
X_19167__328 clknet_1_0__leaf__02748_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__inv_2
X_18446__85 clknet_1_0__leaf__02439_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__inv_2
XFILLER_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19737_ clknet_leaf_91_i_clk _00668_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_16949_ _09553_ _09554_ vssd1 vssd1 vccd1 vccd1 _09555_ sky130_fd_sc_hd__nor2_1
XFILLER_38_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19668_ clknet_leaf_11_i_clk _00599_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f3 sky130_fd_sc_hd__dfxtp_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18619_ net53 rbzero.pov.sclk_buffer\[0\] _03337_ vssd1 vssd1 vccd1 vccd1 _02529_
+ sky130_fd_sc_hd__mux2_1
X_19599_ clknet_leaf_45_i_clk _00530_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20512_ clknet_leaf_78_i_clk _01443_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20443_ net503 _01374_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_51_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_146_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20374_ net434 _01305_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_66_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10960_ _03721_ _03725_ _03735_ _03685_ _03745_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__o311a_1
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10891_ _03635_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__buf_6
XFILLER_70_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12630_ _05258_ _05324_ _05386_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__o21ai_1
XFILLER_71_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12561_ _05277_ _05260_ _05317_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__o21bai_1
XFILLER_180_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11512_ rbzero.tex_g1\[37\] rbzero.tex_g1\[36\] _03727_ vssd1 vssd1 vccd1 vccd1 _04295_
+ sky130_fd_sc_hd__mux2_1
X_14300_ rbzero.debug_overlay.playerX\[-3\] _06961_ vssd1 vssd1 vccd1 vccd1 _06988_
+ sky130_fd_sc_hd__nand2_1
X_15280_ _07964_ _07965_ vssd1 vssd1 vccd1 vccd1 _07966_ sky130_fd_sc_hd__nand2_1
XFILLER_157_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12492_ _05158_ _05248_ _05197_ _05207_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__or4b_1
XFILLER_200_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14231_ _06893_ _06908_ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__or2_1
X_11443_ _03619_ _04226_ _03633_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__o21a_1
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_19_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_109_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14162_ _06850_ vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__buf_4
X_11374_ rbzero.tex_g0\[18\] _03617_ _03611_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__a21o_1
XFILLER_164_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13113_ _05864_ _05869_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__or2_1
X_10325_ _03225_ vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__clkbuf_1
X_14093_ rbzero.wall_tracer.visualWallDist\[7\] _03495_ _06791_ rbzero.wall_tracer.trackDistX\[7\]
+ _03497_ vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__o221a_1
XFILLER_180_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17921_ rbzero.pov.spi_buffer\[15\] rbzero.pov.ready_buffer\[15\] _02153_ vssd1 vssd1
+ vccd1 vccd1 _02160_ sky130_fd_sc_hd__mux2_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _05798_ _05799_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__xnor2_1
X_10256_ _03189_ vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_191_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17852_ rbzero.spi_registers.spi_counter\[1\] rbzero.spi_registers.spi_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__or2_1
X_10187_ rbzero.tex_g0\[40\] rbzero.tex_g0\[39\] _03144_ vssd1 vssd1 vccd1 vccd1 _03153_
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16803_ _09194_ _09304_ vssd1 vssd1 vccd1 vccd1 _09411_ sky130_fd_sc_hd__nor2_1
XFILLER_8_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17783_ _02040_ _02041_ _02049_ vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__o21ai_1
X_14995_ _07660_ _07664_ vssd1 vssd1 vccd1 vccd1 _07683_ sky130_fd_sc_hd__nor2_1
XFILLER_75_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19522_ clknet_leaf_49_i_clk _00468_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16734_ _09336_ _09341_ vssd1 vssd1 vccd1 vccd1 _09342_ sky130_fd_sc_hd__and2b_1
X_13946_ _06696_ vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19453_ clknet_leaf_69_i_clk _00011_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rcp_sel\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16665_ _07992_ _09036_ _09272_ vssd1 vssd1 vccd1 vccd1 _09274_ sky130_fd_sc_hd__o21ai_1
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13877_ _06587_ _06600_ _06588_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__mux2_1
XFILLER_201_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18404_ clknet_1_1__leaf__02433_ vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__buf_1
XFILLER_90_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15616_ _08048_ _08173_ vssd1 vssd1 vccd1 vccd1 _08300_ sky130_fd_sc_hd__nand2_1
X_19384_ rbzero.traced_texa\[8\] rbzero.texV\[8\] _02856_ vssd1 vssd1 vccd1 vccd1
+ _02861_ sky130_fd_sc_hd__a21o_1
X_12828_ _05540_ _05543_ _05584_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__o21ai_2
X_16596_ _09129_ _09098_ vssd1 vssd1 vccd1 vccd1 _09205_ sky130_fd_sc_hd__or2b_1
XFILLER_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18335_ rbzero.spi_registers.new_vshift\[1\] rbzero.spi_registers.spi_buffer\[1\]
+ _02401_ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__mux2_1
X_15547_ _07494_ _07138_ _08000_ _08229_ vssd1 vssd1 vccd1 vccd1 _08231_ sky130_fd_sc_hd__o22ai_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12759_ _05515_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__buf_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18266_ _02364_ vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__clkbuf_1
X_15478_ _08032_ _08034_ vssd1 vssd1 vccd1 vccd1 _08163_ sky130_fd_sc_hd__nor2_1
XFILLER_30_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17217_ _01547_ _01549_ _01548_ vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__o21bai_1
X_14429_ _06906_ rbzero.wall_tracer.stepDistX\[-1\] _07114_ _07116_ vssd1 vssd1 vccd1
+ vccd1 _07117_ sky130_fd_sc_hd__a22oi_4
X_18197_ rbzero.floor_leak\[5\] _02311_ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__or2_1
XFILLER_190_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17148_ _01489_ _01491_ vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09970_ _03038_ vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_157_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17079_ _09578_ _09588_ _09586_ vssd1 vssd1 vccd1 vccd1 _09684_ sky130_fd_sc_hd__a21o_1
Xclkbuf_1_1__f__02737_ clknet_0__02737_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02737_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20090_ clknet_leaf_8_i_clk _01021_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_130_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19241__16 clknet_1_0__leaf__02754_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__inv_2
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19221__377 clknet_1_0__leaf__02753_ vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__inv_2
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20426_ net486 _01357_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20357_ net417 _01288_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10110_ _03112_ vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11090_ gpout0.vpos\[6\] _03873_ _03874_ _03460_ _03875_ vssd1 vssd1 vccd1 vccd1
+ _03876_ sky130_fd_sc_hd__a221o_1
X_20288_ net348 _01219_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19115__282 clknet_1_0__leaf__02742_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__inv_2
X_10041_ _03076_ vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18425__66 clknet_1_0__leaf__02437_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__inv_2
XFILLER_57_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13800_ _06436_ _06473_ _06556_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__and3_1
XFILLER_57_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11992_ _03911_ _04732_ _04725_ _04765_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__a31o_1
X_14780_ _07444_ _07467_ vssd1 vssd1 vccd1 vccd1 _07468_ sky130_fd_sc_hd__xor2_1
XFILLER_91_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10943_ _03696_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__buf_4
X_13731_ _05805_ _05995_ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__nor2_1
XFILLER_182_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16450_ _09030_ _09060_ vssd1 vssd1 vccd1 vccd1 _09061_ sky130_fd_sc_hd__xnor2_1
X_10874_ _03659_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__clkbuf_4
X_13662_ _06402_ _06417_ _06418_ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__o21bai_1
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _08084_ _08085_ vssd1 vssd1 vccd1 vccd1 _08086_ sky130_fd_sc_hd__nor2_1
X_12613_ _05356_ _05364_ _05368_ _05369_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__a211o_1
X_16381_ _08888_ _08889_ _08887_ _08886_ vssd1 vssd1 vccd1 vccd1 _08992_ sky130_fd_sc_hd__o31ai_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13593_ _06296_ _06344_ _06349_ vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__a21oi_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18120_ _03872_ _02263_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__nand2_1
X_15332_ _08015_ _08016_ _08017_ vssd1 vssd1 vccd1 vccd1 _08018_ sky130_fd_sc_hd__a21o_4
X_12544_ _05120_ _05234_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__nor2_4
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18051_ _02229_ vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__clkbuf_1
X_15263_ _07943_ _07948_ vssd1 vssd1 vccd1 vccd1 _07949_ sky130_fd_sc_hd__xor2_1
X_12475_ _05228_ _05231_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__nand2_1
XFILLER_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17002_ _09606_ _09607_ vssd1 vssd1 vccd1 vccd1 _09608_ sky130_fd_sc_hd__xor2_1
XFILLER_184_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11426_ rbzero.tex_g0\[37\] rbzero.tex_g0\[36\] _03699_ vssd1 vssd1 vccd1 vccd1 _04210_
+ sky130_fd_sc_hd__mux2_1
XFILLER_126_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14214_ _03490_ rbzero.wall_tracer.stepDistY\[-3\] _04947_ vssd1 vssd1 vccd1 vccd1
+ _06902_ sky130_fd_sc_hd__a21o_1
X_15194_ _07530_ _07138_ _07732_ vssd1 vssd1 vccd1 vccd1 _07881_ sky130_fd_sc_hd__or3_1
XANTENNA_6 _04388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14145_ _06837_ vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__clkbuf_1
X_11357_ rbzero.debug_overlay.playerY\[3\] _04059_ _04138_ _04141_ vssd1 vssd1 vccd1
+ vccd1 _04142_ sky130_fd_sc_hd__a211o_1
XFILLER_180_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10308_ _03216_ vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14076_ rbzero.wall_tracer.trackDistY\[-2\] _06786_ _06801_ vssd1 vssd1 vccd1 vccd1
+ _00437_ sky130_fd_sc_hd__o21a_1
X_11288_ _03474_ _04062_ _04060_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__or3_1
X_17904_ rbzero.pov.spi_buffer\[7\] rbzero.pov.ready_buffer\[7\] _02143_ vssd1 vssd1
+ vccd1 vccd1 _02151_ sky130_fd_sc_hd__mux2_1
X_13027_ _05777_ _05778_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__nand2_1
X_10239_ _03180_ vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18884_ _02259_ _02702_ _02710_ _02279_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__and4b_1
XFILLER_94_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17835_ _02088_ _02092_ _02089_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__a21bo_1
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17766_ _02032_ _02033_ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__xor2_1
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14978_ _07653_ _07659_ _07665_ vssd1 vssd1 vccd1 vccd1 _07666_ sky130_fd_sc_hd__o21ba_1
XFILLER_82_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19505_ clknet_leaf_54_i_clk _00451_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
X_16717_ _08888_ _07961_ vssd1 vssd1 vccd1 vccd1 _09325_ sky130_fd_sc_hd__nor2_1
X_13929_ _05347_ _06643_ _06637_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__o21a_1
X_17697_ rbzero.wall_tracer.rayAddendX\[-1\] _08447_ _01969_ _01714_ vssd1 vssd1 vccd1
+ vccd1 _01970_ sky130_fd_sc_hd__a22o_1
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19436_ _02334_ _02887_ _02888_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__and3_1
XFILLER_90_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16648_ _08108_ _09256_ vssd1 vssd1 vccd1 vccd1 _09257_ sky130_fd_sc_hd__nor2_1
XFILLER_34_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19367_ _02839_ _02840_ _02841_ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__o21ai_1
XFILLER_37_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16579_ _08970_ _09188_ vssd1 vssd1 vccd1 vccd1 _09189_ sky130_fd_sc_hd__nand2_1
XFILLER_176_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18318_ _02393_ vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19298_ _02785_ _02786_ _02788_ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__or3_1
XFILLER_175_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18249_ rbzero.spi_registers.new_vshift\[3\] _02348_ _02353_ _02314_ vssd1 vssd1
+ vccd1 vccd1 _00798_ sky130_fd_sc_hd__o211a_1
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20211_ net271 _01142_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20142_ clknet_leaf_12_i_clk _01073_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[0\] sky130_fd_sc_hd__dfxtp_2
X_09953_ rbzero.tex_r0\[23\] rbzero.tex_r0\[22\] _03028_ vssd1 vssd1 vccd1 vccd1 _03030_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20073_ clknet_leaf_84_i_clk _01004_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-1\]
+ sky130_fd_sc_hd__dfxtp_4
X_09884_ _02993_ vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__clkbuf_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10590_ rbzero.wall_tracer.visualWallDist\[-1\] rbzero.wall_tracer.visualWallDist\[-2\]
+ rbzero.wall_tracer.visualWallDist\[-3\] _03385_ vssd1 vssd1 vccd1 vccd1 _03386_
+ sky130_fd_sc_hd__or4_1
XFILLER_51_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12260_ rbzero.wall_tracer.mapY\[8\] _04923_ _05017_ vssd1 vssd1 vccd1 vccd1 _05019_
+ sky130_fd_sc_hd__a21o_1
XFILLER_182_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11211_ _03539_ rbzero.row_render.wall\[1\] vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__or2_1
X_20409_ net469 _01340_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12191_ rbzero.wall_tracer.trackDistY\[10\] vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__inv_2
XFILLER_162_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11142_ rbzero.tex_r1\[49\] _03919_ _03926_ _03669_ vssd1 vssd1 vccd1 vccd1 _03927_
+ sky130_fd_sc_hd__a31o_1
XFILLER_107_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 o_gpout[0] sky130_fd_sc_hd__clkbuf_1
XFILLER_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 o_rgb[23] sky130_fd_sc_hd__buf_2
X_11073_ _03854_ rbzero.map_overlay.i_mapdy\[0\] _03856_ rbzero.map_overlay.i_mapdy\[4\]
+ _03858_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__o221a_1
X_15950_ _08562_ _08566_ _08567_ _08522_ vssd1 vssd1 vccd1 vccd1 _08568_ sky130_fd_sc_hd__a31o_1
XFILLER_110_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10024_ rbzero.tex_g1\[52\] rbzero.tex_g1\[53\] _03061_ vssd1 vssd1 vccd1 vccd1 _03067_
+ sky130_fd_sc_hd__mux2_1
X_14901_ _07006_ _07148_ vssd1 vssd1 vccd1 vccd1 _07589_ sky130_fd_sc_hd__or2_1
XFILLER_23_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15881_ _04951_ _03484_ _03458_ _06784_ vssd1 vssd1 vccd1 vccd1 _08506_ sky130_fd_sc_hd__and4b_4
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17620_ rbzero.debug_overlay.playerY\[2\] _01900_ _09620_ vssd1 vssd1 vccd1 vccd1
+ _01901_ sky130_fd_sc_hd__mux2_1
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14832_ _07499_ _07516_ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__nor2_1
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ _01838_ _01839_ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__xnor2_1
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14763_ _06899_ _07177_ vssd1 vssd1 vccd1 vccd1 _07451_ sky130_fd_sc_hd__nor2_1
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ _04743_ _04745_ _04747_ _04748_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__a211o_2
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _08885_ _09008_ _09010_ _09012_ vssd1 vssd1 vccd1 vccd1 _09112_ sky130_fd_sc_hd__a22o_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13714_ _06435_ _06470_ _06426_ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__a21oi_1
X_10926_ rbzero.tex_r0\[29\] rbzero.tex_r0\[28\] _03690_ vssd1 vssd1 vccd1 vccd1 _03712_
+ sky130_fd_sc_hd__mux2_1
X_17482_ _01772_ _01773_ _01774_ _01759_ vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__a211o_1
XFILLER_189_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14694_ _07296_ _07344_ _07347_ _07346_ vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16433_ _09042_ _09043_ vssd1 vssd1 vccd1 vccd1 _09044_ sky130_fd_sc_hd__and2_1
XFILLER_189_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10857_ _03642_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__inv_2
X_13645_ _06392_ _06394_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16364_ _07865_ _08191_ vssd1 vssd1 vccd1 vccd1 _08975_ sky130_fd_sc_hd__nor2_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13576_ _06281_ _06285_ _06332_ vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__a21bo_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ rbzero.traced_texVinit\[8\] rbzero.spi_registers.vshift\[5\] vssd1 vssd1
+ vccd1 vccd1 _03574_ sky130_fd_sc_hd__nand2_1
XFILLER_185_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _02256_ vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__clkbuf_1
X_15315_ _06997_ _08000_ vssd1 vssd1 vccd1 vccd1 _08001_ sky130_fd_sc_hd__nor2_1
XFILLER_9_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12527_ _05277_ _05260_ _05278_ _05283_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__o211a_1
X_16295_ _08905_ _08906_ vssd1 vssd1 vccd1 vccd1 _08907_ sky130_fd_sc_hd__nand2_1
XFILLER_185_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18034_ rbzero.pov.spi_buffer\[69\] rbzero.pov.ready_buffer\[69\] _02142_ vssd1 vssd1
+ vccd1 vccd1 _02219_ sky130_fd_sc_hd__mux2_1
X_15246_ _07931_ _07932_ vssd1 vssd1 vccd1 vccd1 _07933_ sky130_fd_sc_hd__nand2_1
X_12458_ _05213_ _05214_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__xor2_2
X_11409_ rbzero.tex_g0\[49\] rbzero.tex_g0\[48\] _04189_ vssd1 vssd1 vccd1 vccd1 _04193_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15177_ _07862_ _07863_ vssd1 vssd1 vccd1 vccd1 _07864_ sky130_fd_sc_hd__xor2_1
XFILLER_119_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12389_ _03488_ _05143_ _05145_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__a21oi_4
XFILLER_126_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14128_ rbzero.wall_tracer.stepDistX\[1\] _06738_ _06825_ vssd1 vssd1 vccd1 vccd1
+ _06829_ sky130_fd_sc_hd__mux2_1
X_19985_ clknet_leaf_95_i_clk _00916_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14059_ rbzero.wall_tracer.visualWallDist\[-9\] _03496_ _06791_ rbzero.wall_tracer.trackDistX\[-9\]
+ _03485_ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__o221a_1
XFILLER_141_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__02436_ clknet_0__02436_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02436_
+ sky130_fd_sc_hd__clkbuf_16
X_18867_ _02695_ _02696_ _02698_ _02285_ vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__o211a_1
XFILLER_28_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17818_ _01972_ rbzero.debug_overlay.vplaneX\[-1\] _02001_ vssd1 vssd1 vccd1 vccd1
+ _02082_ sky130_fd_sc_hd__a21oi_1
XFILLER_95_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18798_ rbzero.debug_overlay.facingY\[-4\] _02638_ vssd1 vssd1 vccd1 vccd1 _02659_
+ sky130_fd_sc_hd__or2_1
XFILLER_48_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17749_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.debug_overlay.vplaneX\[-6\] _02016_
+ _02017_ vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__and4bb_1
XFILLER_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19419_ _01703_ _01711_ _01710_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__a21oi_1
XFILLER_165_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20125_ clknet_leaf_91_i_clk _01056_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-1\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09936_ rbzero.tex_r0\[31\] rbzero.tex_r0\[30\] _03017_ vssd1 vssd1 vccd1 vccd1 _03021_
+ sky130_fd_sc_hd__mux2_1
XFILLER_132_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20056_ clknet_leaf_7_i_clk _00987_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09867_ net47 rbzero.tex_r0\[63\] _02984_ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__mux2_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09798_ rbzero.tex_r1\[30\] rbzero.tex_r1\[31\] _02943_ vssd1 vssd1 vccd1 vccd1 _02947_
+ sky130_fd_sc_hd__mux2_1
XFILLER_100_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19227__383 clknet_1_1__leaf__02753_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__inv_2
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _03911_ _04515_ _04513_ _04534_ _04537_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__a311o_1
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ gpout0.hpos\[1\] vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__inv_2
XFILLER_199_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _03534_ _03848_ _04390_ _03522_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__a31o_1
XFILLER_201_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13430_ _06118_ _06137_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__xnor2_1
X_10642_ rbzero.map_overlay.i_othery\[1\] _03358_ vssd1 vssd1 vccd1 vccd1 _03438_
+ sky130_fd_sc_hd__xor2_1
XFILLER_186_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13361_ _06078_ _06117_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__and2_1
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10573_ rbzero.map_rom.f1 vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__clkbuf_4
XFILLER_194_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15100_ _07269_ _07333_ _07787_ _07011_ vssd1 vssd1 vccd1 vccd1 _07788_ sky130_fd_sc_hd__o22a_1
XFILLER_181_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12312_ _03480_ _04884_ _04885_ _05068_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__a31o_1
X_16080_ _08407_ _08409_ vssd1 vssd1 vccd1 vccd1 _08694_ sky130_fd_sc_hd__nor2_1
XFILLER_155_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13292_ _05914_ _05915_ _06048_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__a21boi_1
XFILLER_158_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15031_ _06979_ _07281_ _07275_ _07274_ vssd1 vssd1 vccd1 vccd1 _07719_ sky130_fd_sc_hd__o31a_1
XFILLER_5_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12243_ _03495_ _05004_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__nand2_1
XFILLER_142_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12174_ _03374_ _04928_ _04935_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__o21ai_1
XFILLER_123_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11125_ _03504_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__clkbuf_8
X_19770_ clknet_leaf_6_i_clk _00701_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_16982_ _09586_ _09587_ vssd1 vssd1 vccd1 vccd1 _09588_ sky130_fd_sc_hd__nor2_1
XFILLER_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18721_ net61 _02605_ vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__nor2_1
X_11056_ gpout0.vpos\[6\] _03347_ _03363_ _03460_ _03841_ vssd1 vssd1 vccd1 vccd1
+ _03842_ sky130_fd_sc_hd__a221o_1
X_15933_ rbzero.wall_tracer.trackDistX\[-6\] _08508_ _08546_ _08552_ vssd1 vssd1 vccd1
+ vccd1 _00543_ sky130_fd_sc_hd__o22a_1
XFILLER_110_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10007_ rbzero.tex_g1\[60\] rbzero.tex_g1\[61\] _02976_ vssd1 vssd1 vccd1 vccd1 _03058_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18652_ rbzero.pov.ready_buffer\[65\] _06989_ _02539_ vssd1 vssd1 vccd1 vccd1 _02553_
+ sky130_fd_sc_hd__mux2_1
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ rbzero.wall_tracer.mapX\[7\] _08489_ _08488_ _08492_ vssd1 vssd1 vccd1 vccd1
+ _00534_ sky130_fd_sc_hd__a22o_1
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17603_ rbzero.wall_tracer.rayAddendY\[9\] _00013_ _08464_ _01885_ _01887_ vssd1
+ vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__o221a_1
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14815_ _07449_ _07452_ vssd1 vssd1 vccd1 vccd1 _07503_ sky130_fd_sc_hd__xnor2_1
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18583_ rbzero.pov.spi_buffer\[59\] rbzero.pov.spi_buffer\[60\] _02510_ vssd1 vssd1
+ vccd1 vccd1 _02511_ sky130_fd_sc_hd__mux2_1
XFILLER_91_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_100 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_100/HI zeros[9] sky130_fd_sc_hd__conb_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15795_ rbzero.row_render.size\[9\] _08456_ _06738_ _08455_ vssd1 vssd1 vccd1 vccd1
+ _00501_ sky130_fd_sc_hd__a22o_1
Xtop_ew_algofoogle_111 vssd1 vssd1 vccd1 vccd1 ones[4] top_ew_algofoogle_111/LO sky130_fd_sc_hd__conb_1
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_122 vssd1 vssd1 vccd1 vccd1 ones[15] top_ew_algofoogle_122/LO sky130_fd_sc_hd__conb_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17534_ _01805_ _01823_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__xnor2_1
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14746_ _06871_ _06993_ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__nor2_1
X_11958_ net28 net27 vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__and2_1
XFILLER_178_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10909_ rbzero.tex_r0\[17\] rbzero.tex_r0\[16\] _03649_ vssd1 vssd1 vccd1 vccd1 _03695_
+ sky130_fd_sc_hd__mux2_1
X_17465_ _01757_ rbzero.wall_tracer.rayAddendY\[0\] vssd1 vssd1 vccd1 vccd1 _01759_
+ sky130_fd_sc_hd__and2_1
XFILLER_199_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14677_ _07363_ _07364_ vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__nor2_1
X_11889_ _04621_ _04644_ _04663_ _04664_ vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__o31a_2
XFILLER_60_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16416_ _08917_ _08920_ _09026_ vssd1 vssd1 vccd1 vccd1 _09027_ sky130_fd_sc_hd__a21o_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13628_ _05697_ _06056_ _06384_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__nand3_1
X_17396_ _08471_ _08480_ _08469_ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__a21oi_1
XFILLER_158_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16347_ _08524_ _08958_ vssd1 vssd1 vccd1 vccd1 _08959_ sky130_fd_sc_hd__and2_1
XFILLER_9_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13559_ _06121_ _06122_ _05987_ _06035_ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__or4_1
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16278_ _08888_ _08889_ vssd1 vssd1 vccd1 vccd1 _08890_ sky130_fd_sc_hd__nor2_1
XFILLER_172_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18017_ _02210_ vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15229_ _07914_ _07915_ vssd1 vssd1 vccd1 vccd1 _07916_ sky130_fd_sc_hd__nor2_1
XFILLER_201_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19968_ net197 _00899_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09721_ gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__inv_2
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19899_ clknet_leaf_16_i_clk _00830_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_83_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20108_ clknet_leaf_77_i_clk _01039_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
X_09919_ rbzero.tex_r0\[39\] rbzero.tex_r0\[38\] _03006_ vssd1 vssd1 vccd1 vccd1 _03012_
+ sky130_fd_sc_hd__mux2_1
XFILLER_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12930_ _05646_ _05686_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__xnor2_1
X_20039_ clknet_leaf_6_i_clk _00970_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _05609_ _05551_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__nor2_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _07239_ _07263_ _07286_ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__nand3_1
XFILLER_27_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _03782_ _04568_ _04570_ _03865_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__a22o_1
X_15580_ _08262_ _08263_ vssd1 vssd1 vccd1 vccd1 _08264_ sky130_fd_sc_hd__xnor2_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12792_ _05494_ _05488_ _05489_ _05495_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__o31ai_4
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18395__38 clknet_1_0__leaf__02435_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__inv_2
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _07212_ _07218_ vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ net50 _04512_ _04520_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__a21o_1
XFILLER_199_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ rbzero.wall_tracer.trackDistY\[-2\] _01558_ _01583_ _08577_ vssd1 vssd1 vccd1
+ vccd1 _00569_ sky130_fd_sc_hd__o22a_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _06850_ _05064_ vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__nand2_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11674_ rbzero.tex_b1\[15\] rbzero.tex_b1\[14\] _03615_ vssd1 vssd1 vccd1 vccd1 _04455_
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16201_ _08812_ _08813_ vssd1 vssd1 vccd1 vccd1 _08814_ sky130_fd_sc_hd__xor2_1
X_13413_ _05538_ _06098_ _06169_ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__a21o_1
XFILLER_155_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10625_ rbzero.map_overlay.i_mapdx\[3\] rbzero.map_overlay.i_mapdx\[2\] rbzero.map_overlay.i_mapdx\[1\]
+ rbzero.map_overlay.i_mapdx\[0\] vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__or4_1
X_17181_ rbzero.wall_tracer.trackDistY\[-11\] rbzero.wall_tracer.stepDistY\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__nand2_1
XFILLER_167_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14393_ _06900_ _06968_ vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__nor2_1
XFILLER_183_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__02439_ clknet_0__02439_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02439_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_139_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16132_ _07735_ _07786_ _08339_ vssd1 vssd1 vccd1 vccd1 _08745_ sky130_fd_sc_hd__or3_1
XFILLER_6_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13344_ _06090_ _06092_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__xor2_1
X_10556_ rbzero.map_rom.d6 vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__clkinv_2
XFILLER_155_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16063_ _03493_ rbzero.wall_tracer.stepDistY\[9\] _04950_ vssd1 vssd1 vccd1 vccd1
+ _08677_ sky130_fd_sc_hd__a21oi_1
X_10487_ rbzero.tex_b0\[25\] rbzero.tex_b0\[24\] _03302_ vssd1 vssd1 vccd1 vccd1 _03310_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13275_ _05978_ _06031_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__xor2_4
XFILLER_136_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15014_ _07372_ _07701_ vssd1 vssd1 vccd1 vccd1 _07702_ sky130_fd_sc_hd__xnor2_4
X_12226_ _04985_ rbzero.wall_tracer.trackDistX\[-2\] vssd1 vssd1 vccd1 vccd1 _04988_
+ sky130_fd_sc_hd__or2_1
XFILLER_155_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12157_ _04918_ _04878_ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__nor2_1
X_19822_ clknet_leaf_14_i_clk _00753_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11108_ gpout0.vpos\[0\] _03890_ rbzero.debug_overlay.playerX\[-1\] _03783_ _03893_
+ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__a221o_1
XFILLER_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16965_ _09325_ _09433_ vssd1 vssd1 vccd1 vccd1 _09571_ sky130_fd_sc_hd__nand2_1
X_19753_ clknet_leaf_94_i_clk _00684_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_12088_ rbzero.debug_overlay.facingY\[-5\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__and2_1
XFILLER_96_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11039_ rbzero.floor_leak\[2\] _03606_ _03823_ rbzero.floor_leak\[1\] _03824_ vssd1
+ vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__a221o_1
X_18704_ rbzero.debug_overlay.playerY\[-7\] _02588_ _02593_ _02586_ vssd1 vssd1 vccd1
+ vccd1 _01013_ sky130_fd_sc_hd__o211a_1
X_15916_ _08512_ _08536_ _08537_ _08522_ vssd1 vssd1 vccd1 vccd1 _08538_ sky130_fd_sc_hd__a31o_1
X_19684_ clknet_leaf_70_i_clk _00615_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16896_ _09501_ _09502_ vssd1 vssd1 vccd1 vccd1 _09503_ sky130_fd_sc_hd__nor2_1
XFILLER_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18635_ rbzero.pov.ready_buffer\[60\] _06912_ _02540_ vssd1 vssd1 vccd1 vccd1 _02541_
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15847_ _08475_ _08476_ vssd1 vssd1 vccd1 vccd1 _08477_ sky130_fd_sc_hd__and2_1
XFILLER_92_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18566_ rbzero.pov.spi_buffer\[51\] rbzero.pov.spi_buffer\[52\] _02499_ vssd1 vssd1
+ vccd1 vccd1 _02502_ sky130_fd_sc_hd__mux2_1
XFILLER_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ _03474_ _04019_ _04053_ _03911_ vssd1 vssd1 vccd1 vccd1 _08450_ sky130_fd_sc_hd__and4_2
XFILLER_45_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17517_ _04109_ rbzero.debug_overlay.vplaneY\[-6\] _01807_ vssd1 vssd1 vccd1 vccd1
+ _01808_ sky130_fd_sc_hd__or3_1
X_14729_ _07070_ _07071_ vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__or2_1
X_18497_ _02465_ vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__clkbuf_1
XFILLER_162_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17448_ _01722_ _01742_ _01743_ _08460_ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__a31o_1
XFILLER_123_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17379_ _03342_ _09620_ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__nor2_1
XFILLER_119_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20390_ net450 _01321_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19144__307 clknet_1_1__leaf__02746_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__inv_2
XFILLER_55_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10410_ rbzero.tex_b0\[62\] rbzero.tex_b0\[61\] _03269_ vssd1 vssd1 vccd1 vccd1 _03270_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11390_ _04172_ _04173_ _03635_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__mux2_1
XFILLER_165_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19038__212 clknet_1_1__leaf__02735_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__inv_2
XFILLER_125_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10341_ rbzero.tex_b1\[30\] rbzero.tex_b1\[31\] _03232_ vssd1 vssd1 vccd1 vccd1 _03234_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19190__349 clknet_1_1__leaf__02750_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__inv_2
XFILLER_139_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13060_ _05814_ _05816_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__nand2_1
X_10272_ _03197_ vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12011_ _04779_ net62 vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__or2_1
XFILLER_79_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16750_ _09007_ _09142_ _09256_ _09009_ vssd1 vssd1 vccd1 vccd1 _09358_ sky130_fd_sc_hd__o22ai_1
XFILLER_171_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13962_ _06675_ _06709_ _06710_ vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__a21oi_2
XFILLER_101_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15701_ _08249_ _08383_ vssd1 vssd1 vccd1 vccd1 _08384_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12913_ _05667_ _05668_ _05669_ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__a21oi_1
X_16681_ _09172_ _09173_ vssd1 vssd1 vccd1 vccd1 _09290_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13893_ _05265_ _05271_ _06636_ _06648_ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__a31o_1
X_19084__254 clknet_1_0__leaf__02739_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__inv_2
X_15632_ rbzero.wall_tracer.visualWallDist\[10\] _07256_ vssd1 vssd1 vccd1 vccd1 _08315_
+ sky130_fd_sc_hd__nand2_2
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _05529_ _05531_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__xor2_1
XFILLER_61_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _02410_ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__clkbuf_4
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _07581_ vssd1 vssd1 vccd1 vccd1 _08247_ sky130_fd_sc_hd__buf_2
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _05529_ _05531_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__and2b_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ rbzero.wall_tracer.trackDistY\[6\] rbzero.wall_tracer.stepDistY\[6\] vssd1
+ vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__nor2_1
XFILLER_199_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _07193_ _07197_ _07201_ vssd1 vssd1 vccd1 vccd1 _07202_ sky130_fd_sc_hd__o21a_1
X_18282_ _02373_ vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__clkbuf_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _04503_ _04487_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__nor2_1
XFILLER_30_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _08177_ _08178_ vssd1 vssd1 vccd1 vccd1 _08179_ sky130_fd_sc_hd__or2_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17233_ _01566_ _01567_ _01568_ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__a21oi_1
XFILLER_147_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14445_ _04831_ _07132_ _06985_ vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__o21ai_1
X_11657_ rbzero.tex_b1\[27\] _03696_ _03697_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__and3_1
XFILLER_156_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17164_ _09696_ _01507_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__xnor2_1
XFILLER_122_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10608_ _03345_ rbzero.map_rom.a6 rbzero.map_rom.i_row\[4\] _03392_ vssd1 vssd1 vccd1
+ vccd1 _03404_ sky130_fd_sc_hd__or4_1
XFILLER_70_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14376_ _07010_ _07063_ vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__xnor2_1
X_11588_ rbzero.tex_b0\[14\] _03617_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__and2_1
XFILLER_183_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16115_ _08615_ _08631_ _08629_ vssd1 vssd1 vccd1 vccd1 _08728_ sky130_fd_sc_hd__a21o_1
XFILLER_128_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13327_ _05990_ _06074_ _05988_ _06082_ _06083_ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__o32a_1
XFILLER_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17095_ _09630_ _09604_ _09699_ vssd1 vssd1 vccd1 vccd1 _09700_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_1_1__f__02753_ clknet_0__02753_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02753_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10539_ rbzero.vga_sync.vsync vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__inv_6
XFILLER_7_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16046_ _08637_ _08659_ vssd1 vssd1 vccd1 vccd1 _08660_ sky130_fd_sc_hd__xnor2_2
XFILLER_115_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13258_ _05609_ _05990_ _05472_ _05491_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__or4b_1
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12209_ rbzero.wall_tracer.trackDistY\[-5\] vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__inv_2
XFILLER_124_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13189_ _05896_ _05894_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__nor2_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19805_ clknet_leaf_2_i_clk _00736_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17997_ rbzero.pov.spi_buffer\[51\] rbzero.pov.ready_buffer\[51\] _02197_ vssd1 vssd1
+ vccd1 vccd1 _02200_ sky130_fd_sc_hd__mux2_1
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16948_ _09488_ _09489_ _09486_ vssd1 vssd1 vccd1 vccd1 _09554_ sky130_fd_sc_hd__a21oi_1
X_19736_ clknet_leaf_92_i_clk _00667_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16879_ _09014_ _09036_ _09485_ vssd1 vssd1 vccd1 vccd1 _09486_ sky130_fd_sc_hd__nor3_1
XFILLER_37_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19667_ clknet_leaf_11_i_clk _00598_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f4 sky130_fd_sc_hd__dfxtp_1
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18618_ _02528_ vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19598_ clknet_leaf_44_i_clk _00529_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18549_ rbzero.pov.spi_buffer\[43\] rbzero.pov.spi_buffer\[44\] _02488_ vssd1 vssd1
+ vccd1 vccd1 _02493_ sky130_fd_sc_hd__mux2_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20511_ clknet_leaf_78_i_clk _01442_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20442_ net502 _01373_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20373_ net433 _01304_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18452__89 clknet_1_0__leaf__02441_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__inv_2
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10890_ rbzero.tex_r0\[11\] rbzero.tex_r0\[10\] _03663_ vssd1 vssd1 vccd1 vccd1 _03676_
+ sky130_fd_sc_hd__mux2_1
XFILLER_110_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12560_ _05198_ _05225_ _05252_ _05287_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__o211a_1
XFILLER_196_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11511_ rbzero.tex_g1\[38\] _03733_ _03660_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__a21o_1
XFILLER_129_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12491_ _05189_ _05225_ _05231_ _05192_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__or4b_1
X_14230_ _06908_ _06917_ vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__nor2_1
XFILLER_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11442_ _03936_ _03630_ _03639_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__nor3_1
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18912__98 clknet_1_1__leaf__02723_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__inv_2
X_11373_ rbzero.tex_g0\[19\] _04155_ _04156_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__and3_1
X_14161_ _06849_ vssd1 vssd1 vccd1 vccd1 _06850_ sky130_fd_sc_hd__clkbuf_4
XFILLER_180_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10324_ rbzero.tex_b1\[38\] rbzero.tex_b1\[39\] _03221_ vssd1 vssd1 vccd1 vccd1 _03225_
+ sky130_fd_sc_hd__mux2_1
X_13112_ _05867_ _05868_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__xor2_1
X_14092_ rbzero.wall_tracer.trackDistX\[6\] _06788_ _06809_ vssd1 vssd1 vccd1 vccd1
+ _00445_ sky130_fd_sc_hd__o21a_1
XFILLER_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10255_ rbzero.tex_g0\[8\] rbzero.tex_g0\[7\] _03188_ vssd1 vssd1 vccd1 vccd1 _03189_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17920_ _02159_ vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__clkbuf_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ _05798_ _05799_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__or2b_1
XFILLER_26_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17851_ rbzero.spi_registers.spi_counter\[1\] rbzero.spi_registers.spi_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__and2_1
XFILLER_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10186_ _03152_ vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16802_ _09408_ _09409_ vssd1 vssd1 vccd1 vccd1 _09410_ sky130_fd_sc_hd__nand2_1
XFILLER_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17782_ rbzero.wall_tracer.rayAddendX\[5\] _08460_ _02048_ _03497_ vssd1 vssd1 vccd1
+ vccd1 _02049_ sky130_fd_sc_hd__o2bb2a_1
X_14994_ _07647_ _07675_ _07681_ _07676_ vssd1 vssd1 vccd1 vccd1 _07682_ sky130_fd_sc_hd__o211a_1
XFILLER_78_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16733_ _09339_ _09340_ vssd1 vssd1 vccd1 vccd1 _09341_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19521_ clknet_leaf_50_i_clk _00467_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_13945_ rbzero.wall_tracer.stepDistY\[-5\] _06695_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _06696_ sky130_fd_sc_hd__mux2_1
X_18949__132 clknet_1_1__leaf__02726_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__inv_2
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19452_ _02898_ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__clkbuf_1
X_16664_ _07992_ _08391_ _09272_ vssd1 vssd1 vccd1 vccd1 _09273_ sky130_fd_sc_hd__or3_1
XFILLER_35_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13876_ _06632_ vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15615_ _08297_ _08298_ vssd1 vssd1 vccd1 vccd1 _08299_ sky130_fd_sc_hd__and2_2
XFILLER_62_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19383_ rbzero.traced_texa\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _02860_
+ sky130_fd_sc_hd__nand2_1
X_12827_ _05544_ _05554_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__or2_1
X_16595_ _09186_ _09187_ vssd1 vssd1 vccd1 vccd1 _09204_ sky130_fd_sc_hd__or2_1
XFILLER_62_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18334_ _02402_ vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__clkbuf_1
X_15546_ _08229_ _07138_ _08102_ vssd1 vssd1 vccd1 vccd1 _08230_ sky130_fd_sc_hd__or3_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _05376_ _05390_ _05514_ _05416_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__o31a_4
XFILLER_61_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11709_ net3 vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__buf_2
X_18265_ rbzero.spi_registers.spi_buffer\[2\] rbzero.spi_registers.new_sky\[2\] _02361_
+ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__mux2_1
X_15477_ _08115_ _08161_ vssd1 vssd1 vccd1 vccd1 _08162_ sky130_fd_sc_hd__xnor2_2
X_12689_ _05414_ _05359_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__or2_1
XFILLER_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17216_ rbzero.wall_tracer.trackDistY\[-6\] rbzero.wall_tracer.stepDistY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__nand2_1
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14428_ _03491_ _07115_ _06906_ vssd1 vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__a21oi_1
X_18196_ rbzero.spi_registers.new_leak\[4\] _02310_ _02317_ _02314_ vssd1 vssd1 vccd1
+ vccd1 _00781_ sky130_fd_sc_hd__o211a_1
XFILLER_144_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17147_ _01490_ _09648_ _09646_ vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__a21oi_1
X_14359_ _04839_ rbzero.wall_tracer.stepDistX\[-9\] _07043_ _07046_ vssd1 vssd1 vccd1
+ vccd1 _07047_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_183_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18995__174 clknet_1_0__leaf__02730_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__inv_2
XFILLER_115_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17078_ _09681_ _09682_ vssd1 vssd1 vccd1 vccd1 _09683_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_1__f__02736_ clknet_0__02736_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02736_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16029_ _07735_ vssd1 vssd1 vccd1 vccd1 _08643_ sky130_fd_sc_hd__buf_2
XFILLER_171_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19719_ clknet_leaf_95_i_clk _00650_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20425_ net485 _01356_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20356_ net416 _01287_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20287_ net347 _01218_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ rbzero.tex_g1\[45\] rbzero.tex_g1\[46\] _03073_ vssd1 vssd1 vccd1 vccd1 _03076_
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11991_ net44 _04731_ _04725_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__and3_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13730_ _05536_ _06155_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__nor2_1
X_10942_ rbzero.tex_r0\[41\] rbzero.tex_r0\[40\] _03727_ vssd1 vssd1 vccd1 vccd1 _03728_
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13661_ _06403_ _06404_ _06416_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__and3_1
X_10873_ _03610_ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__buf_4
XFILLER_72_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15400_ _08076_ _07976_ _08083_ vssd1 vssd1 vccd1 vccd1 _08085_ sky130_fd_sc_hd__and3_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _05224_ _05226_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__nor2_4
X_16380_ _08989_ _08990_ vssd1 vssd1 vccd1 vccd1 _08991_ sky130_fd_sc_hd__xor2_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _06345_ _06348_ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__nor2_1
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15331_ _04841_ rbzero.wall_tracer.stepDistX\[7\] vssd1 vssd1 vccd1 vccd1 _08017_
+ sky130_fd_sc_hd__nor2_1
XFILLER_196_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12543_ _05274_ _05285_ _05299_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__or3_2
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19122__287 clknet_1_0__leaf__02744_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__inv_2
XFILLER_184_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19196__355 clknet_1_0__leaf__02750_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__inv_2
XFILLER_157_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18050_ rbzero.spi_registers.spi_buffer\[1\] rbzero.spi_registers.spi_buffer\[0\]
+ _02227_ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__mux2_1
X_15262_ _07946_ _07947_ vssd1 vssd1 vccd1 vccd1 _07948_ sky130_fd_sc_hd__xor2_1
X_12474_ _05229_ _05230_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__xor2_2
XFILLER_8_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17001_ _09428_ _09506_ _09505_ vssd1 vssd1 vccd1 vccd1 _09607_ sky130_fd_sc_hd__a21boi_1
XFILLER_144_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14213_ _06893_ _06900_ vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__nor2_1
X_11425_ _04207_ _04208_ _03739_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__mux2_1
XFILLER_184_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15193_ _07581_ _07138_ vssd1 vssd1 vccd1 vccd1 _07880_ sky130_fd_sc_hd__nor2_1
XFILLER_137_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_7 _04828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14144_ rbzero.wall_tracer.stepDistX\[9\] _06779_ _04833_ vssd1 vssd1 vccd1 vccd1
+ _06837_ sky130_fd_sc_hd__mux2_1
XFILLER_126_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11356_ rbzero.debug_overlay.playerY\[4\] _04064_ _04092_ rbzero.debug_overlay.playerY\[-3\]
+ _04140_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__a221o_1
XFILLER_153_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10307_ rbzero.tex_b1\[46\] rbzero.tex_b1\[47\] _03210_ vssd1 vssd1 vccd1 vccd1 _03216_
+ sky130_fd_sc_hd__mux2_1
X_14075_ rbzero.wall_tracer.visualWallDist\[-2\] _06796_ _06791_ rbzero.wall_tracer.trackDistX\[-2\]
+ _06797_ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__o221a_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11287_ _04070_ _04071_ _04055_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__a21bo_1
XFILLER_106_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17903_ _02150_ vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__clkbuf_1
X_13026_ _05771_ _05772_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__xor2_1
X_10238_ rbzero.tex_g0\[16\] rbzero.tex_g0\[15\] _03177_ vssd1 vssd1 vccd1 vccd1 _03180_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18883_ _04507_ _04500_ _04499_ _04508_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__a31o_1
XFILLER_117_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19016__192 clknet_1_1__leaf__02733_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__inv_2
XFILLER_94_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10169_ _02982_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__buf_4
X_17834_ rbzero.wall_tracer.rayAddendX\[9\] _03509_ _08464_ _02093_ _02096_ vssd1
+ vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__o221a_1
XFILLER_48_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14977_ _07660_ _07664_ vssd1 vssd1 vccd1 vccd1 _07665_ sky130_fd_sc_hd__and2_1
X_17765_ _02012_ _02014_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__or2b_1
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19504_ clknet_leaf_54_i_clk _00450_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_50_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16716_ _08643_ _08191_ vssd1 vssd1 vccd1 vccd1 _09324_ sky130_fd_sc_hd__nor2_1
X_13928_ _06680_ vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__clkbuf_1
X_17696_ _04100_ _01968_ vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__xor2_1
XFILLER_63_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16647_ _08134_ vssd1 vssd1 vccd1 vccd1 _09256_ sky130_fd_sc_hd__buf_2
X_19435_ gpout1.clk_div\[0\] gpout1.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__or2_1
XFILLER_62_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13859_ _06565_ _06564_ vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__and2b_1
XFILLER_23_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16578_ _09186_ _09187_ vssd1 vssd1 vccd1 vccd1 _09188_ sky130_fd_sc_hd__xor2_1
X_19366_ _02844_ _02845_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__nand2_1
XFILLER_124_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15529_ _08211_ _08212_ vssd1 vssd1 vccd1 vccd1 _08213_ sky130_fd_sc_hd__nor2_1
X_18317_ rbzero.spi_registers.new_other\[4\] rbzero.spi_registers.spi_buffer\[4\]
+ _02388_ vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__mux2_1
X_19297_ rbzero.traced_texa\[-6\] rbzero.texV\[-6\] _02787_ vssd1 vssd1 vccd1 vccd1
+ _02788_ sky130_fd_sc_hd__o21ai_1
XFILLER_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18248_ rbzero.spi_registers.vshift\[3\] _02349_ vssd1 vssd1 vccd1 vccd1 _02353_
+ sky130_fd_sc_hd__or2_1
XFILLER_124_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18179_ rbzero.spi_registers.new_mapd\[3\] _02289_ _02307_ _02301_ vssd1 vssd1 vccd1
+ vccd1 _00774_ sky130_fd_sc_hd__o211a_1
XFILLER_117_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20210_ net270 _01141_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20141_ clknet_leaf_32_i_clk _01072_ vssd1 vssd1 vccd1 vccd1 rbzero.hsync sky130_fd_sc_hd__dfxtp_2
X_09952_ _03029_ vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20072_ clknet_leaf_83_i_clk _01003_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-2\]
+ sky130_fd_sc_hd__dfxtp_4
X_09883_ rbzero.tex_r0\[56\] rbzero.tex_r0\[55\] _02984_ vssd1 vssd1 vccd1 vccd1 _02993_
+ sky130_fd_sc_hd__mux2_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_18_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18430__70 clknet_1_0__leaf__02438_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__inv_2
XFILLER_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11210_ _03967_ _03976_ _03985_ _03994_ _03718_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__o221a_1
X_20408_ net468 _01339_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[63\] sky130_fd_sc_hd__dfxtp_1
X_12190_ _03483_ _03458_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__nand2_1
XFILLER_179_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11141_ _03620_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__clkbuf_4
X_20339_ net399 _01270_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[58\] sky130_fd_sc_hd__dfxtp_1
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 o_gpout[1] sky130_fd_sc_hd__clkbuf_1
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 o_rgb[6] sky130_fd_sc_hd__buf_2
XFILLER_1_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11072_ _03854_ rbzero.map_overlay.i_mapdy\[0\] rbzero.map_overlay.i_mapdy\[3\] _03857_
+ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_163_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10023_ _03066_ vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14900_ _07556_ _07587_ vssd1 vssd1 vccd1 vccd1 _07588_ sky130_fd_sc_hd__nand2_2
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15880_ _08488_ _08504_ _08505_ _08489_ rbzero.wall_tracer.mapX\[10\] vssd1 vssd1
+ vccd1 vccd1 _00537_ sky130_fd_sc_hd__a32o_1
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14831_ _07497_ _07518_ vssd1 vssd1 vccd1 vccd1 _07519_ sky130_fd_sc_hd__nor2_1
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ _01811_ _01820_ _01821_ _01805_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__a22o_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14762_ _06899_ _07156_ vssd1 vssd1 vccd1 vccd1 _07450_ sky130_fd_sc_hd__or2_1
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ clknet_1_0__leaf__04486_ _04730_ _04725_ _04726_ vssd1 vssd1 vccd1 vccd1
+ _04748_ sky130_fd_sc_hd__a31o_2
XFILLER_56_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16501_ _08643_ _09110_ _08989_ _08988_ vssd1 vssd1 vccd1 vccd1 _09111_ sky130_fd_sc_hd__o31ai_1
XFILLER_45_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13713_ _06436_ _06469_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__and2_1
X_10925_ rbzero.tex_r0\[31\] _03696_ _03697_ _03659_ vssd1 vssd1 vccd1 vccd1 _03711_
+ sky130_fd_sc_hd__a31o_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17481_ _01757_ rbzero.wall_tracer.rayAddendY\[0\] _01756_ vssd1 vssd1 vccd1 vccd1
+ _01774_ sky130_fd_sc_hd__o21a_1
X_14693_ _07377_ _07380_ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__xnor2_1
XFILLER_189_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__02739_ clknet_0__02739_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02739_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19220_ clknet_1_0__leaf__02743_ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__buf_1
X_16432_ _09032_ _09033_ _09041_ vssd1 vssd1 vccd1 vccd1 _09043_ sky130_fd_sc_hd__nand3_1
XFILLER_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13644_ _06376_ _06375_ _06359_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__a21o_1
X_10856_ rbzero.row_render.side _03641_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__nor2_1
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19204__362 clknet_1_1__leaf__02751_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__inv_2
XFILLER_198_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _08907_ _08883_ vssd1 vssd1 vccd1 vccd1 _08974_ sky130_fd_sc_hd__or2b_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13575_ _06330_ _06331_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__nand2_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10787_ rbzero.traced_texVinit\[8\] rbzero.spi_registers.vshift\[5\] vssd1 vssd1
+ vccd1 vccd1 _03573_ sky130_fd_sc_hd__or2_1
X_18102_ rbzero.spi_registers.sclk_buffer\[2\] rbzero.spi_registers.sclk_buffer\[1\]
+ _04834_ vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__mux2_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15314_ _07141_ vssd1 vssd1 vccd1 vccd1 _08000_ sky130_fd_sc_hd__clkbuf_4
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12526_ _05221_ _05182_ _05224_ _05282_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__o22a_1
XFILLER_184_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16294_ _08794_ _08884_ _08904_ vssd1 vssd1 vccd1 vccd1 _08906_ sky130_fd_sc_hd__nand3_1
XFILLER_158_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18033_ _02218_ vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15245_ _07929_ _07930_ vssd1 vssd1 vccd1 vccd1 _07932_ sky130_fd_sc_hd__or2_1
X_12457_ _05105_ _05127_ _05131_ _05199_ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__o31a_1
XFILLER_138_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11408_ _03656_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__buf_4
XFILLER_158_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15176_ _07084_ _07281_ vssd1 vssd1 vccd1 vccd1 _07863_ sky130_fd_sc_hd__nor2_1
X_12388_ _05067_ _04873_ _04887_ _05144_ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__o31a_1
XFILLER_99_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14127_ _06828_ vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__clkbuf_1
X_11339_ _04116_ _04123_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__or2_1
XFILLER_193_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19984_ clknet_leaf_0_i_clk _00915_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14058_ _05005_ vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__clkbuf_4
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13009_ _05760_ _05765_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1__f__02435_ clknet_0__02435_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02435_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_95_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18866_ _02258_ _02694_ _02697_ rbzero.vga_sync.vsync vssd1 vssd1 vccd1 vccd1 _02698_
+ sky130_fd_sc_hd__a31o_1
XFILLER_121_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17817_ _01972_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__inv_2
X_18797_ rbzero.pov.ready_buffer\[26\] _02644_ _02658_ _02651_ vssd1 vssd1 vccd1 vccd1
+ _01041_ sky130_fd_sc_hd__a211o_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17748_ rbzero.debug_overlay.vplaneX\[-1\] _04100_ vssd1 vssd1 vccd1 vccd1 _02017_
+ sky130_fd_sc_hd__nand2_1
XFILLER_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17679_ rbzero.debug_overlay.vplaneX\[-3\] rbzero.wall_tracer.rayAddendX\[-3\] vssd1
+ vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__nand2_1
XFILLER_36_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19418_ rbzero.wall_tracer.rayAddendY\[-7\] _02868_ _08454_ _02877_ vssd1 vssd1 vccd1
+ vccd1 _01443_ sky130_fd_sc_hd__a22o_1
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19349_ _02831_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__inv_2
XFILLER_176_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20124_ clknet_leaf_90_i_clk _01055_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-2\]
+ sky130_fd_sc_hd__dfxtp_4
X_09935_ _03020_ vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20055_ clknet_leaf_87_i_clk _00986_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[71\]
+ sky130_fd_sc_hd__dfxtp_1
X_09866_ _02983_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__clkbuf_4
XFILLER_131_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09797_ _02946_ vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__clkbuf_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10710_ _03493_ _03496_ _03498_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__o21a_1
XFILLER_159_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _03896_ _04470_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__and2_1
XFILLER_198_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10641_ rbzero.map_overlay.i_othery\[0\] vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__inv_2
XFILLER_158_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13360_ _06076_ _06077_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__or2_1
XFILLER_194_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10572_ _03349_ _03356_ _03367_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__or3_1
XFILLER_194_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12311_ rbzero.wall_tracer.visualWallDist\[2\] _05067_ _03488_ vssd1 vssd1 vccd1
+ vccd1 _05068_ sky130_fd_sc_hd__a21o_1
X_13291_ _06023_ _06040_ _06047_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__or3_1
XFILLER_108_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15030_ _07716_ _07717_ vssd1 vssd1 vccd1 vccd1 _07718_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12242_ rbzero.wall_tracer.trackDistX\[10\] _04953_ _04955_ _05003_ vssd1 vssd1 vccd1
+ vccd1 _05004_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_181_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12173_ _03390_ _04934_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__nand2_1
XFILLER_150_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11124_ _03906_ _03908_ _03909_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__a21o_4
XFILLER_96_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16981_ _09580_ _09585_ vssd1 vssd1 vccd1 vccd1 _09587_ sky130_fd_sc_hd__nor2_1
XFILLER_7_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18720_ _07016_ _02604_ _02587_ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__mux2_1
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11055_ _03840_ rbzero.debug_overlay.playerY\[4\] rbzero.debug_overlay.playerX\[2\]
+ _03782_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__a22o_1
X_15932_ _08550_ _08551_ _08507_ vssd1 vssd1 vccd1 vccd1 _08552_ sky130_fd_sc_hd__o21ai_1
XFILLER_114_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10006_ _03057_ vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18651_ _02534_ _02551_ _02552_ _02356_ vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__o211a_1
X_15863_ _08490_ _08491_ vssd1 vssd1 vccd1 vccd1 _08492_ sky130_fd_sc_hd__xnor2_1
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17602_ _01872_ _01875_ _01886_ _03497_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__a211o_1
X_14814_ _07501_ _07485_ vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__xnor2_1
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18582_ _02442_ vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__buf_4
X_15794_ rbzero.row_render.size\[8\] _08456_ _06733_ _08455_ vssd1 vssd1 vccd1 vccd1
+ _00500_ sky130_fd_sc_hd__a22o_1
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_101 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_101/HI zeros[10]
+ sky130_fd_sc_hd__conb_1
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_112 vssd1 vssd1 vccd1 vccd1 ones[5] top_ew_algofoogle_112/LO sky130_fd_sc_hd__conb_1
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ _01821_ _01822_ vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__and2_1
X_14745_ _07428_ _07432_ vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__or2b_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ net28 net27 vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__and2b_1
XFILLER_91_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19128__293 clknet_1_1__leaf__02744_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__inv_2
X_10908_ _03691_ _03692_ _03693_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__mux2_1
X_17464_ _01757_ rbzero.wall_tracer.rayAddendY\[0\] vssd1 vssd1 vccd1 vccd1 _01758_
+ sky130_fd_sc_hd__nor2_1
X_14676_ _07340_ _07362_ vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__and2_1
XFILLER_189_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11888_ _04314_ _04622_ _04623_ _04632_ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__nand4_1
XFILLER_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16415_ _09013_ _09025_ vssd1 vssd1 vccd1 vccd1 _09026_ sky130_fd_sc_hd__xnor2_1
X_13627_ _05862_ _05995_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__nor2_1
XFILLER_60_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10839_ rbzero.row_render.texu\[4\] rbzero.row_render.texu\[3\] vssd1 vssd1 vccd1
+ vccd1 _03625_ sky130_fd_sc_hd__nand2_1
XFILLER_60_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17395_ _01695_ vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16346_ _08954_ _08957_ vssd1 vssd1 vccd1 vccd1 _08958_ sky130_fd_sc_hd__xnor2_4
X_13558_ _06121_ _05988_ _06061_ _06122_ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__o22ai_2
X_19065_ clknet_1_0__leaf__02732_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__buf_1
XFILLER_145_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12509_ _05252_ _05255_ _05260_ _05264_ _05265_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__a41o_1
X_16277_ _07857_ vssd1 vssd1 vccd1 vccd1 _08889_ sky130_fd_sc_hd__clkbuf_4
X_13489_ _06008_ _06071_ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__nor2_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15228_ _07727_ _07774_ _07773_ vssd1 vssd1 vccd1 vccd1 _07915_ sky130_fd_sc_hd__a21oi_1
X_18016_ rbzero.pov.spi_buffer\[60\] rbzero.pov.ready_buffer\[60\] _02208_ vssd1 vssd1
+ vccd1 vccd1 _02210_ sky130_fd_sc_hd__mux2_1
XFILLER_173_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15159_ _07844_ _07845_ vssd1 vssd1 vccd1 vccd1 _07846_ sky130_fd_sc_hd__xnor2_1
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19967_ net196 _00898_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09720_ gpout0.hpos\[8\] vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__clkbuf_4
XFILLER_132_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19898_ clknet_leaf_16_i_clk _00829_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18849_ rbzero.debug_overlay.vplaneY\[-3\] _02660_ vssd1 vssd1 vccd1 vccd1 _02687_
+ sky130_fd_sc_hd__or2_1
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09918_ _03011_ vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__clkbuf_1
X_20107_ clknet_leaf_77_i_clk _01038_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_19_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20038_ clknet_leaf_6_i_clk _00969_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[54\]
+ sky130_fd_sc_hd__dfxtp_1
X_09849_ _02973_ vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ _05494_ _05616_ _05595_ _05591_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__a31o_1
XFILLER_2_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _04586_ _04587_ net18 vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__mux2_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12791_ _05392_ _05496_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__nor2_1
XFILLER_61_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _07141_ _07213_ _07216_ _07217_ vssd1 vssd1 vccd1 vccd1 _07218_ sky130_fd_sc_hd__o31a_1
XFILLER_26_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ net51 _04519_ _04516_ net53 vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__a22o_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _06746_ _07130_ vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__xnor2_1
X_11673_ rbzero.tex_b1\[13\] rbzero.tex_b1\[12\] _03616_ vssd1 vssd1 vccd1 vccd1 _04454_
+ sky130_fd_sc_hd__mux2_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16200_ _08671_ _08691_ _08690_ vssd1 vssd1 vccd1 vccd1 _08813_ sky130_fd_sc_hd__a21oi_2
XFILLER_30_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13412_ _06123_ _06128_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__nand2_1
XFILLER_128_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17180_ _01522_ vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__clkbuf_4
X_10624_ rbzero.map_overlay.i_mapdx\[4\] vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__inv_2
XFILLER_168_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14392_ _07078_ _06970_ vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_0__f__02438_ clknet_0__02438_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02438_
+ sky130_fd_sc_hd__clkbuf_16
X_16131_ _07735_ _07332_ vssd1 vssd1 vccd1 vccd1 _08744_ sky130_fd_sc_hd__nor2_1
XFILLER_139_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13343_ _05549_ _06098_ _06099_ _06097_ vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__a211o_1
XFILLER_139_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10555_ rbzero.wall_tracer.mapY\[5\] vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__inv_2
XFILLER_6_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16062_ _08672_ _08675_ vssd1 vssd1 vccd1 vccd1 _08676_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13274_ _06029_ _06030_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__and2_1
X_10486_ _03309_ vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15013_ _07471_ _07476_ _07475_ vssd1 vssd1 vccd1 vccd1 _07701_ sky130_fd_sc_hd__a21o_1
X_12225_ _04985_ rbzero.wall_tracer.trackDistX\[-2\] rbzero.wall_tracer.trackDistX\[-3\]
+ _04986_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__a22o_1
XFILLER_123_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19821_ clknet_leaf_14_i_clk _00752_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12156_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[9\] vssd1
+ vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__nor2_1
XFILLER_155_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11107_ rbzero.debug_overlay.playerX\[-2\] _03527_ vssd1 vssd1 vccd1 vccd1 _03893_
+ sky130_fd_sc_hd__xor2_1
X_19752_ clknet_leaf_90_i_clk _00683_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_16964_ _09568_ _09569_ vssd1 vssd1 vccd1 vccd1 _09570_ sky130_fd_sc_hd__xor2_1
X_12087_ _04845_ _04848_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__or2_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18703_ rbzero.pov.ready_buffer\[46\] _02413_ _02582_ _02592_ vssd1 vssd1 vccd1 vccd1
+ _02593_ sky130_fd_sc_hd__a211o_1
X_11038_ rbzero.floor_leak\[1\] _03610_ _03662_ rbzero.floor_leak\[0\] vssd1 vssd1
+ vccd1 vccd1 _03824_ sky130_fd_sc_hd__o211a_1
X_15915_ _08533_ _08534_ _08535_ vssd1 vssd1 vccd1 vccd1 _08537_ sky130_fd_sc_hd__a21o_1
X_19683_ clknet_leaf_70_i_clk _00614_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16895_ _09388_ _09391_ _09500_ vssd1 vssd1 vccd1 vccd1 _09502_ sky130_fd_sc_hd__and3_1
XFILLER_92_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18634_ _02539_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__clkbuf_4
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ _03353_ _06914_ vssd1 vssd1 vccd1 vccd1 _08476_ sky130_fd_sc_hd__or2_1
XFILLER_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18565_ _02501_ vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__clkbuf_1
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12989_ _05733_ _05745_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__xnor2_1
X_15777_ _08448_ vssd1 vssd1 vccd1 vccd1 _08449_ sky130_fd_sc_hd__buf_4
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17516_ _01805_ _01806_ vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__nand2_1
X_14728_ _07400_ _07402_ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__nand2_1
X_19061__233 clknet_1_1__leaf__02737_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__inv_2
X_18496_ rbzero.pov.spi_buffer\[18\] rbzero.pov.spi_buffer\[19\] _02455_ vssd1 vssd1
+ vccd1 vccd1 _02465_ sky130_fd_sc_hd__mux2_1
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17447_ rbzero.debug_overlay.vplaneY\[-6\] _01732_ vssd1 vssd1 vccd1 vccd1 _01743_
+ sky130_fd_sc_hd__or2_1
XFILLER_60_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14659_ _07091_ _07177_ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__nor2_1
XFILLER_159_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17378_ _03395_ _08472_ vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__or2_1
XFILLER_186_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16329_ _08938_ _08939_ vssd1 vssd1 vccd1 vccd1 _08941_ sky130_fd_sc_hd__and2_1
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10340_ _03233_ vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_191_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10271_ rbzero.tex_b1\[63\] net49 _03117_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__mux2_1
XFILLER_3_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12010_ _04779_ _04314_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__nand2_1
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13961_ _06675_ _06677_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__nor2_1
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15700_ _08381_ _08382_ vssd1 vssd1 vccd1 vccd1 _08383_ sky130_fd_sc_hd__nor2_1
XFILLER_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12912_ _05392_ _05465_ _05534_ _05538_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__and4b_1
X_16680_ _09267_ _09288_ vssd1 vssd1 vccd1 vccd1 _09289_ sky130_fd_sc_hd__xnor2_2
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13892_ _06637_ _06647_ _06630_ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__a21o_1
XFILLER_34_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15631_ _08190_ _08219_ _08313_ vssd1 vssd1 vccd1 vccd1 _08314_ sky130_fd_sc_hd__a21boi_1
X_12843_ _05574_ _05599_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__xor2_1
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15562_ _08245_ _07766_ vssd1 vssd1 vccd1 vccd1 _08246_ sky130_fd_sc_hd__nor2_1
X_18350_ net40 net39 vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__or2_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _05524_ _05530_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__nor2_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _07198_ _07199_ _07200_ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__or3_1
X_17301_ rbzero.wall_tracer.trackDistY\[5\] _01558_ _01627_ _09308_ vssd1 vssd1 vccd1
+ vccd1 _00576_ sky130_fd_sc_hd__o22a_1
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _03834_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__clkbuf_4
X_18281_ rbzero.spi_registers.spi_buffer\[2\] rbzero.spi_registers.new_floor\[2\]
+ _02370_ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__mux2_1
X_15493_ _08054_ _08057_ _08176_ vssd1 vssd1 vccd1 vccd1 _08178_ sky130_fd_sc_hd__and3_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14444_ _04920_ _05075_ _06850_ vssd1 vssd1 vccd1 vccd1 _07132_ sky130_fd_sc_hd__mux2_1
X_17232_ _01560_ _01562_ _01561_ vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__o21bai_1
XFILLER_175_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11656_ rbzero.tex_b1\[25\] rbzero.tex_b1\[24\] _04376_ vssd1 vssd1 vccd1 vccd1 _04437_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17163_ _01477_ _01506_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__xnor2_1
X_10607_ _03353_ _03345_ _03400_ _03402_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__a211o_1
XFILLER_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14375_ _07015_ _07062_ vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11587_ _04366_ _04367_ _04368_ _03740_ _03702_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__o221a_1
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16114_ _08725_ _08726_ vssd1 vssd1 vccd1 vccd1 _08727_ sky130_fd_sc_hd__nor2_1
XFILLER_116_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13326_ _05990_ _05988_ _06061_ _05472_ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__o22a_1
X_17094_ _09693_ _09698_ vssd1 vssd1 vccd1 vccd1 _09699_ sky130_fd_sc_hd__xor2_1
XFILLER_183_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__02752_ clknet_0__02752_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02752_
+ sky130_fd_sc_hd__clkbuf_16
X_10538_ _03336_ vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16045_ _08657_ _08658_ vssd1 vssd1 vccd1 vccd1 _08659_ sky130_fd_sc_hd__nand2_1
XFILLER_127_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13257_ _05491_ _05696_ _05472_ _05609_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__o2bb2a_1
X_10469_ _03300_ vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12208_ rbzero.wall_tracer.trackDistY\[-4\] vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__inv_2
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13188_ _05891_ _05893_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__nor2_1
XFILLER_151_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19804_ clknet_leaf_3_i_clk _00735_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12139_ _04899_ _04900_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__nand2_1
XFILLER_2_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17996_ _02199_ vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19735_ clknet_leaf_93_i_clk _00666_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16947_ _09551_ _09552_ vssd1 vssd1 vccd1 vccd1 _09553_ sky130_fd_sc_hd__or2_1
XFILLER_81_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19666_ clknet_leaf_4_i_clk _00597_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_16878_ _09016_ _08678_ vssd1 vssd1 vccd1 vccd1 _09485_ sky130_fd_sc_hd__or2_1
XFILLER_37_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18617_ rbzero.pov.ss_buffer\[1\] rbzero.pov.ss_buffer\[0\] _04827_ vssd1 vssd1 vccd1
+ vccd1 _02528_ sky130_fd_sc_hd__mux2_1
X_15829_ rbzero.traced_texa\[8\] _08463_ _08462_ rbzero.wall_tracer.visualWallDist\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__a22o_1
X_19597_ clknet_leaf_44_i_clk _00528_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18926__111 clknet_1_0__leaf__02724_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__inv_2
X_18548_ _02492_ vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18479_ _02456_ vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20510_ clknet_leaf_82_i_clk _01441_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20441_ net501 _01372_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20372_ net432 _01303_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18972__153 clknet_1_0__leaf__02728_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__inv_2
XFILLER_102_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19068__239 clknet_1_0__leaf__02738_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__inv_2
XFILLER_84_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11510_ rbzero.tex_g1\[39\] _03729_ _03730_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__and3_1
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12490_ _05229_ _05230_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__xnor2_2
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11441_ _03538_ _03539_ _03640_ _03996_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__o31ai_1
XFILLER_20_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14160_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__buf_2
X_11372_ _03697_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__clkbuf_4
XFILLER_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13111_ _05609_ _05499_ _05467_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__a21oi_1
X_10323_ _03224_ vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14091_ rbzero.wall_tracer.visualWallDist\[6\] _03495_ _06784_ rbzero.wall_tracer.trackDistY\[6\]
+ _03497_ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__o221a_1
XFILLER_180_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13042_ _05726_ _05759_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__xor2_1
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10254_ _03143_ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__buf_4
XFILLER_65_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17850_ _02107_ rbzero.spi_registers.spi_cmd\[1\] _02110_ vssd1 vssd1 vccd1 vccd1
+ _02111_ sky130_fd_sc_hd__and3_1
X_10185_ rbzero.tex_g0\[41\] rbzero.tex_g0\[40\] _03144_ vssd1 vssd1 vccd1 vccd1 _03152_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16801_ _09405_ _09407_ vssd1 vssd1 vccd1 vccd1 _09409_ sky130_fd_sc_hd__nand2_1
XFILLER_66_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17781_ _02046_ _02047_ vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__xnor2_1
X_14993_ _07647_ _07678_ _07679_ _07623_ _07680_ vssd1 vssd1 vccd1 vccd1 _07681_ sky130_fd_sc_hd__a221o_1
XFILLER_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19520_ clknet_leaf_50_i_clk _00466_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16732_ _08862_ _09110_ vssd1 vssd1 vccd1 vccd1 _09340_ sky130_fd_sc_hd__nor2_1
X_13944_ _06637_ _06688_ _06689_ _06694_ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__a31o_2
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19451_ _04828_ _02896_ _02897_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__and3_1
X_16663_ _09270_ _09271_ vssd1 vssd1 vccd1 vccd1 _09272_ sky130_fd_sc_hd__xnor2_1
X_13875_ rbzero.wall_tracer.stepDistY\[-11\] _06631_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _06632_ sky130_fd_sc_hd__mux2_1
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15614_ _08183_ _08296_ vssd1 vssd1 vccd1 vccd1 _08298_ sky130_fd_sc_hd__or2_1
X_12826_ _05575_ _05582_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__xor2_1
X_19382_ rbzero.traced_texa\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _02859_
+ sky130_fd_sc_hd__or2_1
XFILLER_34_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16594_ rbzero.wall_tracer.trackDistX\[4\] _08553_ _09197_ _09203_ vssd1 vssd1 vccd1
+ vccd1 _00553_ sky130_fd_sc_hd__o22a_1
XFILLER_90_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18333_ rbzero.spi_registers.new_vshift\[0\] rbzero.spi_registers.spi_buffer\[0\]
+ _02401_ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__mux2_1
X_15545_ _07273_ vssd1 vssd1 vccd1 vccd1 _08229_ sky130_fd_sc_hd__buf_2
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _05380_ _05331_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__nand2_1
XFILLER_72_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15476_ _08159_ _08160_ vssd1 vssd1 vccd1 vccd1 _08161_ sky130_fd_sc_hd__nor2_1
X_18264_ _02363_ vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__clkbuf_1
XFILLER_187_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12688_ _05347_ _05363_ _05444_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__a21o_1
X_17215_ rbzero.wall_tracer.trackDistY\[-6\] rbzero.wall_tracer.stepDistY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__or2_1
X_14427_ rbzero.wall_tracer.stepDistY\[-1\] vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__inv_2
X_11639_ rbzero.tex_b1\[59\] _03696_ _03697_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__and3_1
X_18195_ rbzero.floor_leak\[4\] _02311_ vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__or2_1
XFILLER_129_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17146_ _09641_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__inv_2
XFILLER_156_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14358_ _06852_ _06658_ _07045_ _06985_ vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__o211ai_1
X_19173__334 clknet_1_1__leaf__02748_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__inv_2
X_13309_ _06058_ _06064_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__and2_1
X_17077_ _09680_ _09673_ vssd1 vssd1 vccd1 vccd1 _09682_ sky130_fd_sc_hd__and2b_1
Xclkbuf_1_1__f__02735_ clknet_0__02735_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02735_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_144_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14289_ _04838_ rbzero.wall_tracer.stepDistX\[-7\] _06973_ _06976_ vssd1 vssd1 vccd1
+ vccd1 _06977_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16028_ _07735_ _07270_ _08641_ vssd1 vssd1 vccd1 vccd1 _08642_ sky130_fd_sc_hd__or3_1
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17979_ _02190_ vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__clkbuf_1
X_19718_ clknet_leaf_0_i_clk _00649_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19649_ clknet_leaf_45_i_clk _00580_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20424_ net484 _01355_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20355_ net415 _01286_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20286_ net346 _01217_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11990_ net43 _04730_ _04725_ _04726_ net42 vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__a32o_1
XFILLER_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10941_ _03649_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__buf_4
XFILLER_44_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__02755_ clknet_0__02755_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02755_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13660_ _06403_ _06404_ _06416_ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__a21oi_1
X_10872_ _03653_ _03657_ _03607_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__mux2_1
XFILLER_182_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12611_ _05365_ _05366_ _05367_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__mux2_1
XFILLER_71_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _06298_ _06346_ _06347_ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__a21o_1
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _03493_ rbzero.wall_tracer.stepDistY\[7\] _04950_ vssd1 vssd1 vccd1 vccd1
+ _08016_ sky130_fd_sc_hd__a21oi_1
XFILLER_197_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ _05298_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__clkbuf_2
XFILLER_157_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15261_ _06873_ _07839_ vssd1 vssd1 vccd1 vccd1 _07947_ sky130_fd_sc_hd__nor2_1
X_12473_ _05094_ _05132_ _05199_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__o21a_1
XFILLER_8_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17000_ _09604_ _09605_ vssd1 vssd1 vccd1 vccd1 _09606_ sky130_fd_sc_hd__nand2_1
X_18979__159 clknet_1_1__leaf__02729_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__inv_2
XFILLER_126_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14212_ _06899_ vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__clkbuf_4
X_11424_ rbzero.tex_g0\[35\] rbzero.tex_g0\[34\] _04188_ vssd1 vssd1 vccd1 vccd1 _04208_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15192_ _07877_ _07878_ _07744_ _07743_ vssd1 vssd1 vccd1 vccd1 _07879_ sky130_fd_sc_hd__o31ai_2
XFILLER_125_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_8 _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14143_ _06836_ vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__clkbuf_1
X_11355_ rbzero.debug_overlay.playerY\[0\] _04079_ _04081_ rbzero.debug_overlay.playerY\[-9\]
+ _04139_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__a221o_1
XFILLER_125_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10306_ _03215_ vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14074_ rbzero.wall_tracer.trackDistY\[-3\] _06786_ _06800_ vssd1 vssd1 vccd1 vccd1
+ _00436_ sky130_fd_sc_hd__o21a_1
X_11286_ _03460_ _04040_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__nand2_1
XFILLER_152_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17902_ rbzero.pov.spi_buffer\[6\] rbzero.pov.ready_buffer\[6\] _02143_ vssd1 vssd1
+ vccd1 vccd1 _02150_ sky130_fd_sc_hd__mux2_1
X_13025_ _05779_ _05780_ _05781_ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__a21o_1
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10237_ _03179_ vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18882_ _08439_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__buf_4
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17833_ _02082_ _02085_ _02095_ _03497_ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__a211o_1
XFILLER_39_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10168_ _03142_ vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18416__57 clknet_1_1__leaf__02437_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__inv_2
X_17764_ _01985_ rbzero.wall_tracer.rayAddendX\[4\] vssd1 vssd1 vccd1 vccd1 _02032_
+ sky130_fd_sc_hd__xor2_1
XFILLER_82_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10099_ rbzero.tex_g1\[17\] rbzero.tex_g1\[18\] _03106_ vssd1 vssd1 vccd1 vccd1 _03107_
+ sky130_fd_sc_hd__mux2_1
X_14976_ _07648_ _07663_ vssd1 vssd1 vccd1 vccd1 _07664_ sky130_fd_sc_hd__and2_1
X_19503_ clknet_leaf_40_i_clk _00449_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[10\]
+ sky130_fd_sc_hd__dfxtp_4
X_16715_ _09266_ _09246_ vssd1 vssd1 vccd1 vccd1 _09323_ sky130_fd_sc_hd__or2b_1
XFILLER_75_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13927_ rbzero.wall_tracer.stepDistY\[-7\] _06679_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _06680_ sky130_fd_sc_hd__mux2_1
X_17695_ rbzero.debug_overlay.vplaneX\[-6\] rbzero.debug_overlay.vplaneX\[-7\] rbzero.debug_overlay.vplaneX\[-8\]
+ _01967_ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__o31a_1
XFILLER_74_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19434_ gpout1.clk_div\[0\] gpout1.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__nand2_1
X_16646_ _09253_ _09254_ vssd1 vssd1 vccd1 vccd1 _09255_ sky130_fd_sc_hd__nand2_1
X_13858_ _05324_ _06614_ vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__nor2_1
XFILLER_62_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19365_ rbzero.traced_texa\[6\] rbzero.texV\[6\] vssd1 vssd1 vccd1 vccd1 _02845_
+ sky130_fd_sc_hd__nand2_1
X_12809_ _05561_ _05564_ _05565_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__a21oi_1
XFILLER_37_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16577_ _08972_ _09070_ _09068_ vssd1 vssd1 vccd1 vccd1 _09187_ sky130_fd_sc_hd__a21oi_1
X_13789_ _06439_ _06545_ vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__nand2_1
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18316_ _02392_ vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__clkbuf_1
XFILLER_163_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15528_ _08210_ _08203_ vssd1 vssd1 vccd1 vccd1 _08212_ sky130_fd_sc_hd__and2b_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19296_ rbzero.traced_texa\[-6\] rbzero.texV\[-6\] _02783_ vssd1 vssd1 vccd1 vccd1
+ _02787_ sky130_fd_sc_hd__a21o_1
XFILLER_163_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18247_ rbzero.spi_registers.new_vshift\[2\] _02348_ _02352_ _02314_ vssd1 vssd1
+ vccd1 vccd1 _00797_ sky130_fd_sc_hd__o211a_1
X_15459_ _08015_ _08016_ _08017_ vssd1 vssd1 vccd1 vccd1 _08144_ sky130_fd_sc_hd__a21oi_2
XFILLER_191_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18178_ rbzero.mapdxw\[1\] _02291_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__or2_1
XFILLER_184_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17129_ _01466_ _01472_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09951_ rbzero.tex_r0\[24\] rbzero.tex_r0\[23\] _03028_ vssd1 vssd1 vccd1 vccd1 _03029_
+ sky130_fd_sc_hd__mux2_1
XFILLER_144_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20140_ clknet_leaf_26_i_clk _01071_ vssd1 vssd1 vccd1 vccd1 rbzero.vga_sync.vsync
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_0__02749_ _02749_ vssd1 vssd1 vccd1 vccd1 clknet_0__02749_ sky130_fd_sc_hd__clkbuf_16
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09882_ _02992_ vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__clkbuf_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20071_ clknet_leaf_64_i_clk _01002_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-3\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20407_ net467 _01338_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11140_ _03733_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__clkbuf_4
XFILLER_134_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20338_ net398 _01269_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[57\] sky130_fd_sc_hd__dfxtp_1
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 o_gpout[2] sky130_fd_sc_hd__clkbuf_1
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 o_rgb[7] sky130_fd_sc_hd__buf_2
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11071_ gpout0.vpos\[6\] vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__inv_2
X_20269_ net329 _01200_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10022_ rbzero.tex_g1\[53\] rbzero.tex_g1\[54\] _03061_ vssd1 vssd1 vccd1 vccd1 _03066_
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14830_ _07487_ _07493_ _07496_ vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__and3_1
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11973_ gpout4.clk_div\[1\] _04732_ _04725_ _04746_ vssd1 vssd1 vccd1 vccd1 _04747_
+ sky130_fd_sc_hd__a31o_1
XFILLER_45_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14761_ _06939_ _07147_ vssd1 vssd1 vccd1 vccd1 _07449_ sky130_fd_sc_hd__nor2_1
XFILLER_99_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16500_ _08081_ vssd1 vssd1 vccd1 vccd1 _09110_ sky130_fd_sc_hd__clkbuf_4
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10924_ rbzero.tex_r0\[30\] _03709_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__and2_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ _06438_ _06468_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__nor2_1
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17480_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__or2_1
X_14692_ _06901_ _07378_ _07379_ vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__a21bo_1
Xclkbuf_1_0__f__02738_ clknet_0__02738_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02738_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16431_ _09032_ _09033_ _09041_ vssd1 vssd1 vccd1 vccd1 _09042_ sky130_fd_sc_hd__a21o_1
X_10855_ rbzero.row_render.wall\[0\] _03640_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__nand2_1
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13643_ _06376_ _06359_ _06375_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__nand3_1
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16362_ _08860_ _08877_ _08875_ vssd1 vssd1 vccd1 vccd1 _08973_ sky130_fd_sc_hd__a21o_1
XFILLER_169_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13574_ _06228_ _06277_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__xor2_1
X_10786_ _03568_ _03571_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__nand2_1
XFILLER_12_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18101_ _02255_ vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__clkbuf_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15313_ _07996_ _07998_ vssd1 vssd1 vccd1 vccd1 _07999_ sky130_fd_sc_hd__nor2_1
X_12525_ _05197_ _05281_ _05207_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__o21a_1
X_16293_ _08794_ _08884_ _08904_ vssd1 vssd1 vccd1 vccd1 _08905_ sky130_fd_sc_hd__a21o_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18032_ rbzero.pov.spi_buffer\[68\] rbzero.pov.ready_buffer\[68\] _02208_ vssd1 vssd1
+ vccd1 vccd1 _02218_ sky130_fd_sc_hd__mux2_1
X_12456_ _05097_ _05099_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__and2_1
X_15244_ _07929_ _07930_ vssd1 vssd1 vccd1 vccd1 _07931_ sky130_fd_sc_hd__nand2_1
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11407_ _04187_ _04190_ _03740_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__mux2_1
X_15175_ _07713_ _07860_ _07861_ vssd1 vssd1 vccd1 vccd1 _07862_ sky130_fd_sc_hd__a21bo_1
X_12387_ rbzero.wall_tracer.visualWallDist\[-1\] _05067_ _03487_ vssd1 vssd1 vccd1
+ vccd1 _05144_ sky130_fd_sc_hd__a21oi_1
XFILLER_153_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14126_ rbzero.wall_tracer.stepDistX\[0\] _06733_ _06825_ vssd1 vssd1 vccd1 vccd1
+ _06828_ sky130_fd_sc_hd__mux2_1
X_11338_ rbzero.debug_overlay.facingX\[-1\] _04093_ _04122_ vssd1 vssd1 vccd1 vccd1
+ _04123_ sky130_fd_sc_hd__a21oi_1
X_19983_ net212 _00914_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14057_ rbzero.wall_tracer.trackDistX\[-10\] _06788_ _06790_ vssd1 vssd1 vccd1 vccd1
+ _00429_ sky130_fd_sc_hd__o21a_1
XFILLER_193_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11269_ _04053_ _03511_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__nand2b_1
XFILLER_98_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13008_ _05764_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__inv_2
XFILLER_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__02434_ clknet_0__02434_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02434_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_122_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18865_ _04507_ _04499_ _04500_ _04508_ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__and4bb_1
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17816_ _02078_ _02079_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__nor2_1
XFILLER_95_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18796_ rbzero.debug_overlay.facingY\[-5\] _02645_ vssd1 vssd1 vccd1 vccd1 _02658_
+ sky130_fd_sc_hd__and2_1
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17747_ rbzero.debug_overlay.vplaneX\[-1\] _04100_ vssd1 vssd1 vccd1 vccd1 _02016_
+ sky130_fd_sc_hd__or2_1
X_14959_ _06866_ _07646_ vssd1 vssd1 vccd1 vccd1 _07647_ sky130_fd_sc_hd__or2_1
XFILLER_35_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17678_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.wall_tracer.rayAddendX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__and2_1
XFILLER_62_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19417_ _01708_ _02876_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__xnor2_1
X_16629_ _09228_ _09236_ vssd1 vssd1 vccd1 vccd1 _09238_ sky130_fd_sc_hd__nor2_1
XFILLER_165_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19348_ _02828_ _02829_ _02830_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__and3_1
XFILLER_176_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19279_ rbzero.traced_texa\[-8\] rbzero.texV\[-8\] vssd1 vssd1 vccd1 vccd1 _02773_
+ sky130_fd_sc_hd__nand2_1
XFILLER_164_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20123_ clknet_leaf_91_i_clk _01054_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
X_09934_ rbzero.tex_r0\[32\] rbzero.tex_r0\[31\] _03017_ vssd1 vssd1 vccd1 vccd1 _03020_
+ sky130_fd_sc_hd__mux2_1
X_09865_ _02982_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__buf_4
X_20054_ clknet_leaf_87_i_clk _00985_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09796_ rbzero.tex_r1\[31\] rbzero.tex_r1\[32\] _02943_ vssd1 vssd1 vccd1 vccd1 _02946_
+ sky130_fd_sc_hd__mux2_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ rbzero.map_overlay.i_othery\[4\] rbzero.map_rom.i_row\[4\] vssd1 vssd1 vccd1
+ vccd1 _03436_ sky130_fd_sc_hd__xor2_1
XFILLER_186_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10571_ _03357_ _03358_ _03361_ _03366_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__a211o_1
XFILLER_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12310_ _05066_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__buf_2
XFILLER_158_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13290_ _06044_ _06046_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__xnor2_1
XFILLER_177_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12241_ _04955_ _05001_ _05002_ _04953_ rbzero.wall_tracer.trackDistX\[10\] vssd1
+ vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__a32oi_2
XFILLER_170_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12172_ _03358_ _04928_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11123_ gpout0.vpos\[9\] vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__clkbuf_4
XFILLER_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16980_ _09580_ _09585_ vssd1 vssd1 vccd1 vccd1 _09586_ sky130_fd_sc_hd__and2_1
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_64_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11054_ gpout0.vpos\[7\] vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__clkinv_2
X_15931_ _08547_ _08548_ _08549_ _04946_ vssd1 vssd1 vccd1 vccd1 _08551_ sky130_fd_sc_hd__a31o_1
XFILLER_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10005_ rbzero.tex_g1\[61\] rbzero.tex_g1\[62\] _02976_ vssd1 vssd1 vccd1 vccd1 _03057_
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18650_ rbzero.debug_overlay.playerX\[-4\] _02542_ vssd1 vssd1 vccd1 vccd1 _02552_
+ sky130_fd_sc_hd__or2_1
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15862_ rbzero.wall_tracer.mapX\[6\] _07826_ _08483_ vssd1 vssd1 vccd1 vccd1 _08491_
+ sky130_fd_sc_hd__a21boi_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17601_ _01786_ _01757_ _01875_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__o21ba_1
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14813_ _06933_ _07006_ vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__nor2_1
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18581_ _02509_ vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ rbzero.row_render.size\[7\] _08456_ _06726_ _08455_ vssd1 vssd1 vccd1 vccd1
+ _00499_ sky130_fd_sc_hd__a22o_1
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtop_ew_algofoogle_102 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_102/HI zeros[11]
+ sky130_fd_sc_hd__conb_1
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17532_ _01808_ _01811_ _01820_ vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_79_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_91_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_113 vssd1 vssd1 vccd1 vccd1 ones[6] top_ew_algofoogle_113/LO sky130_fd_sc_hd__conb_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14744_ _07429_ _07430_ _07431_ vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__o21ai_1
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ net27 net28 vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__nor2b_2
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10907_ _03635_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__buf_6
X_17463_ rbzero.debug_overlay.vplaneY\[0\] vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__clkbuf_4
X_11887_ _04658_ net14 _04662_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__and3b_1
X_14675_ _07340_ _07362_ vssd1 vssd1 vccd1 vccd1 _07363_ sky130_fd_sc_hd__nor2_1
XFILLER_33_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16414_ _09023_ _09024_ vssd1 vssd1 vccd1 vccd1 _09025_ sky130_fd_sc_hd__nor2_1
X_10838_ _03623_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__buf_6
X_13626_ _05527_ _05995_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__nor2_1
XFILLER_38_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17394_ rbzero.map_rom.i_col\[4\] _01694_ _08506_ vssd1 vssd1 vccd1 vccd1 _01695_
+ sky130_fd_sc_hd__mux2_1
XFILLER_160_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16345_ _08713_ _08715_ _08832_ _08955_ _08956_ vssd1 vssd1 vccd1 vccd1 _08957_ sky130_fd_sc_hd__o311ai_4
XFILLER_9_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18920__106 clknet_1_0__leaf__02723_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__inv_2
X_13557_ _06262_ _06261_ _06173_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__a21o_1
X_10769_ rbzero.traced_texVinit\[2\] rbzero.texV\[2\] _03554_ vssd1 vssd1 vccd1 vccd1
+ _03555_ sky130_fd_sc_hd__o21ai_2
XFILLER_185_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12508_ _05175_ _05182_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__nand2_1
X_16276_ _08000_ vssd1 vssd1 vccd1 vccd1 _08888_ sky130_fd_sc_hd__buf_2
X_13488_ _05503_ _05995_ vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__nor2_1
XFILLER_200_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18015_ _02209_ vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15227_ _07874_ _07913_ vssd1 vssd1 vccd1 vccd1 _07914_ sky130_fd_sc_hd__xnor2_1
X_12439_ _05186_ _05195_ _05153_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_17_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15158_ _07783_ _07789_ _07785_ vssd1 vssd1 vccd1 vccd1 _07845_ sky130_fd_sc_hd__a21oi_1
XFILLER_141_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14109_ rbzero.wall_tracer.stepDistX\[-8\] _06669_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _06819_ sky130_fd_sc_hd__mux2_1
XFILLER_99_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19966_ net195 _00897_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[46\] sky130_fd_sc_hd__dfxtp_1
X_15089_ _07246_ _07290_ _07244_ vssd1 vssd1 vccd1 vccd1 _07777_ sky130_fd_sc_hd__a21oi_1
XFILLER_114_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19897_ clknet_leaf_17_i_clk _00828_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_110_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18848_ rbzero.pov.ready_buffer\[5\] _02666_ _02686_ _02675_ vssd1 vssd1 vccd1 vccd1
+ _01064_ sky130_fd_sc_hd__a211o_1
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18779_ rbzero.debug_overlay.facingX\[-2\] _02638_ vssd1 vssd1 vccd1 vccd1 _02649_
+ sky130_fd_sc_hd__or2_1
XFILLER_94_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20106_ clknet_leaf_77_i_clk _01037_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09917_ rbzero.tex_r0\[40\] rbzero.tex_r0\[39\] _03006_ vssd1 vssd1 vccd1 vccd1 _03011_
+ sky130_fd_sc_hd__mux2_1
XFILLER_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20037_ clknet_leaf_1_i_clk _00968_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_09848_ rbzero.tex_r1\[6\] rbzero.tex_r1\[7\] _02965_ vssd1 vssd1 vccd1 vccd1 _02973_
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ rbzero.tex_r1\[39\] net71 _02932_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__mux2_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ gpout0.hpos\[0\] _03527_ _03526_ _04020_ net15 net16 vssd1 vssd1 vccd1 vccd1
+ _04587_ sky130_fd_sc_hd__mux4_1
XFILLER_160_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12790_ _05493_ _05546_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__nor2_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ net4 net3 vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__and2b_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11672_ _04451_ _04452_ _03739_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__mux2_1
XFILLER_14_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _07147_ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__clkbuf_4
XFILLER_186_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19253__3 clknet_1_0__leaf__02433_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__inv_2
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13411_ _06099_ _06143_ _06167_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__a21oi_1
X_10623_ _03412_ _03418_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__nand2_1
XFILLER_167_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14391_ _07078_ _06968_ vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_0__f__02437_ clknet_0__02437_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02437_
+ sky130_fd_sc_hd__clkbuf_16
X_16130_ _08107_ _07787_ vssd1 vssd1 vccd1 vccd1 _08743_ sky130_fd_sc_hd__nor2_1
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13342_ _05576_ _06055_ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__and2_1
XFILLER_183_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10554_ rbzero.debug_overlay.playerX\[4\] vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__inv_2
XFILLER_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16061_ _08673_ _08674_ vssd1 vssd1 vccd1 vccd1 _08675_ sky130_fd_sc_hd__nand2_1
XFILLER_155_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13273_ _05972_ _06005_ _06028_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__or3_1
X_10485_ rbzero.tex_b0\[26\] rbzero.tex_b0\[25\] _03302_ vssd1 vssd1 vccd1 vccd1 _03309_
+ sky130_fd_sc_hd__mux2_1
XFILLER_154_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12224_ rbzero.wall_tracer.trackDistY\[-3\] vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__inv_2
X_15012_ _07477_ _07526_ _07528_ _07699_ vssd1 vssd1 vccd1 vccd1 _07700_ sky130_fd_sc_hd__a22o_2
XFILLER_154_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19820_ clknet_leaf_14_i_clk _00751_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12155_ _04873_ _04875_ _04876_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__o21a_1
XFILLER_150_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11106_ gpout0.vpos\[0\] _03890_ rbzero.debug_overlay.playerX\[-1\] _03783_ _03891_
+ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__o221a_1
XFILLER_190_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19751_ clknet_leaf_92_i_clk _00682_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16963_ _08888_ _08333_ vssd1 vssd1 vccd1 vccd1 _09569_ sky130_fd_sc_hd__nor2_1
XFILLER_155_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12086_ _04846_ _04847_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__nand2_1
XFILLER_110_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18702_ _06879_ _02535_ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__nor2_1
X_11037_ _03610_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__buf_6
X_15914_ _08533_ _08534_ _08535_ vssd1 vssd1 vccd1 vccd1 _08536_ sky130_fd_sc_hd__nand3_1
X_19682_ clknet_leaf_72_i_clk _00613_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_16894_ _09388_ _09391_ _09500_ vssd1 vssd1 vccd1 vccd1 _09501_ sky130_fd_sc_hd__a21oi_1
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18633_ _02538_ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__clkbuf_4
XFILLER_92_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15845_ _03353_ _07825_ vssd1 vssd1 vccd1 vccd1 _08475_ sky130_fd_sc_hd__nand2_1
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18564_ rbzero.pov.spi_buffer\[50\] rbzero.pov.spi_buffer\[51\] _02499_ vssd1 vssd1
+ vccd1 vccd1 _02501_ sky130_fd_sc_hd__mux2_1
XFILLER_52_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15776_ _08447_ vssd1 vssd1 vccd1 vccd1 _08448_ sky130_fd_sc_hd__buf_4
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _05740_ _05743_ _05744_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a21oi_1
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17515_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.debug_overlay.vplaneY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__nand2_1
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14727_ _07411_ _07414_ vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__nand2_1
X_18495_ _02464_ vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__clkbuf_1
X_11939_ _03537_ _04666_ _04668_ net40 _04713_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__a221o_1
XFILLER_162_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17446_ rbzero.debug_overlay.vplaneY\[-6\] _01732_ vssd1 vssd1 vccd1 vccd1 _01742_
+ sky130_fd_sc_hd__nand2_1
X_14658_ _06787_ _04839_ _06860_ _07114_ vssd1 vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__and4_1
XFILLER_162_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13609_ _06122_ _05991_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__or2_1
X_17377_ _01681_ vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14589_ _06979_ _07052_ vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__nor2_1
XFILLER_146_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16328_ _08938_ _08939_ vssd1 vssd1 vccd1 vccd1 _08940_ sky130_fd_sc_hd__nor2_1
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16259_ _08864_ _08870_ vssd1 vssd1 vccd1 vccd1 _08871_ sky130_fd_sc_hd__and2_1
XFILLER_145_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19949_ net178 _00880_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_6_0_i_clk clknet_2_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_51_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10270_ _03196_ vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13960_ _06690_ _06708_ _06664_ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__mux2_1
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12911_ _05392_ _05526_ _05538_ _05465_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_86_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13891_ _05347_ _06643_ _06645_ _05410_ _06646_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__a221o_1
XFILLER_98_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15630_ _08220_ _08188_ vssd1 vssd1 vccd1 vccd1 _08313_ sky130_fd_sc_hd__or2b_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12842_ _05586_ _05598_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19045__218 clknet_1_0__leaf__02736_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__inv_2
XFILLER_34_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _07530_ vssd1 vssd1 vccd1 vccd1 _08245_ sky130_fd_sc_hd__buf_2
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12773_ _05523_ _05501_ _05512_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__nor3_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _01534_ _01625_ _01626_ _01526_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__a31o_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _07175_ _04948_ _03492_ _07134_ vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__or4_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18280_ _02372_ vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__clkbuf_1
X_11724_ _04496_ _04501_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__nand2_1
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15492_ _08054_ _08057_ _08176_ vssd1 vssd1 vccd1 vccd1 _08177_ sky130_fd_sc_hd__a21oi_1
XFILLER_159_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17231_ rbzero.wall_tracer.trackDistY\[-4\] rbzero.wall_tracer.stepDistY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__nand2_1
X_11655_ _04434_ _04435_ _03739_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__mux2_1
XFILLER_35_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14443_ _07129_ _07130_ vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__nand2_1
XFILLER_122_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17162_ _01494_ _01505_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__xnor2_1
XFILLER_122_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10606_ _03373_ _03352_ rbzero.map_rom.a6 _03401_ rbzero.map_rom.f1 vssd1 vssd1 vccd1
+ vccd1 _03402_ sky130_fd_sc_hd__a2111o_1
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11586_ rbzero.tex_b0\[9\] rbzero.tex_b0\[8\] _03709_ vssd1 vssd1 vccd1 vccd1 _04368_
+ sky130_fd_sc_hd__mux2_1
X_14374_ _07060_ _07061_ vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__and2b_1
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16113_ _08633_ _08722_ _08724_ vssd1 vssd1 vccd1 vccd1 _08726_ sky130_fd_sc_hd__and3_1
XFILLER_128_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10537_ rbzero.tex_b0\[1\] rbzero.tex_b0\[0\] _02983_ vssd1 vssd1 vccd1 vccd1 _03336_
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13325_ _05989_ _06080_ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__nor2_1
X_17093_ _09696_ _09697_ vssd1 vssd1 vccd1 vccd1 _09698_ sky130_fd_sc_hd__and2b_1
Xclkbuf_1_1__f__02751_ clknet_0__02751_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02751_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16044_ _08638_ _08386_ _08656_ vssd1 vssd1 vccd1 vccd1 _08658_ sky130_fd_sc_hd__nand3_1
X_10468_ rbzero.tex_b0\[34\] rbzero.tex_b0\[33\] _03291_ vssd1 vssd1 vccd1 vccd1 _03300_
+ sky130_fd_sc_hd__mux2_1
X_13256_ _06011_ _06012_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__nor2_1
X_12207_ _04965_ _04968_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__nor2_1
X_19238__13 clknet_1_0__leaf__02754_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__inv_2
X_13187_ _05942_ _05943_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__nor2_1
X_10399_ rbzero.tex_b1\[2\] rbzero.tex_b1\[3\] _03254_ vssd1 vssd1 vccd1 vccd1 _03264_
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12138_ _04857_ _04864_ _04852_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__a21o_1
X_19803_ clknet_leaf_3_i_clk _00734_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_17995_ rbzero.pov.spi_buffer\[50\] rbzero.pov.ready_buffer\[50\] _02197_ vssd1 vssd1
+ vccd1 vccd1 _02199_ sky130_fd_sc_hd__mux2_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16946_ _09549_ _09550_ vssd1 vssd1 vccd1 vccd1 _09552_ sky130_fd_sc_hd__nor2_1
X_19734_ clknet_leaf_93_i_clk _00665_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_12069_ _03481_ _03486_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__nor2_1
XFILLER_84_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19665_ clknet_leaf_4_i_clk _00596_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_16877_ _09482_ _09483_ vssd1 vssd1 vccd1 vccd1 _09484_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18616_ _02527_ vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__clkbuf_1
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15828_ rbzero.traced_texa\[7\] _08463_ _08462_ rbzero.wall_tracer.visualWallDist\[7\]
+ vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__a22o_1
X_19596_ clknet_leaf_44_i_clk _00527_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18547_ rbzero.pov.spi_buffer\[42\] rbzero.pov.spi_buffer\[43\] _02488_ vssd1 vssd1
+ vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
X_15759_ _03501_ _03809_ _08439_ vssd1 vssd1 vccd1 vccd1 _08440_ sky130_fd_sc_hd__and3b_1
XFILLER_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18478_ rbzero.pov.spi_buffer\[9\] rbzero.pov.spi_buffer\[10\] _02455_ vssd1 vssd1
+ vccd1 vccd1 _02456_ sky130_fd_sc_hd__mux2_1
XFILLER_166_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17429_ rbzero.debug_overlay.vplaneY\[-3\] rbzero.wall_tracer.rayAddendY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__nor2_1
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20440_ net500 _01371_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20371_ net431 _01302_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19150__313 clknet_1_0__leaf__02746_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__inv_2
XFILLER_173_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11440_ _03688_ _04197_ _04206_ _04223_ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__a31o_1
XFILLER_156_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11371_ _03696_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__clkbuf_4
XFILLER_165_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10322_ rbzero.tex_b1\[39\] rbzero.tex_b1\[40\] _03221_ vssd1 vssd1 vccd1 vccd1 _03224_
+ sky130_fd_sc_hd__mux2_1
X_13110_ _05865_ _05866_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__xnor2_1
X_14090_ rbzero.wall_tracer.trackDistX\[5\] _06788_ _06808_ vssd1 vssd1 vccd1 vccd1
+ _00444_ sky130_fd_sc_hd__o21a_1
XFILLER_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13041_ _05767_ _05797_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__or2_1
XFILLER_106_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10253_ _03187_ vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10184_ _03151_ vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16800_ _09405_ _09407_ vssd1 vssd1 vccd1 vccd1 _09408_ sky130_fd_sc_hd__or2_1
XFILLER_121_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17780_ _02023_ _02026_ _02027_ _02029_ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__o22a_1
X_14992_ _07011_ _07670_ vssd1 vssd1 vccd1 vccd1 _07680_ sky130_fd_sc_hd__or2_1
XFILLER_78_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16731_ _09232_ _09337_ _09338_ vssd1 vssd1 vccd1 vccd1 _09339_ sky130_fd_sc_hd__a21bo_1
XFILLER_115_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13943_ _05476_ _06693_ _06629_ vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__a21o_1
XFILLER_46_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19450_ gpout4.clk_div\[1\] gpout4.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__or2_1
X_16662_ _08247_ _08681_ vssd1 vssd1 vccd1 vccd1 _09271_ sky130_fd_sc_hd__nor2_1
X_13874_ _05210_ _06607_ _06628_ _06630_ vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__a31o_1
XFILLER_74_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15613_ _08183_ _08296_ vssd1 vssd1 vccd1 vccd1 _08297_ sky130_fd_sc_hd__nand2_1
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19381_ _08439_ _02857_ _02858_ _02319_ rbzero.texV\[8\] vssd1 vssd1 vccd1 vccd1
+ _01425_ sky130_fd_sc_hd__a32o_1
X_12825_ _05580_ _05581_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__nand2_1
XFILLER_90_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16593_ _08512_ _09202_ _08489_ vssd1 vssd1 vccd1 vccd1 _09203_ sky130_fd_sc_hd__a21o_1
X_18332_ _02400_ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__clkbuf_4
XFILLER_188_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15544_ _08226_ _08227_ vssd1 vssd1 vccd1 vccd1 _08228_ sky130_fd_sc_hd__xnor2_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12756_ _05505_ _05471_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__or2_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18263_ rbzero.spi_registers.spi_buffer\[1\] rbzero.spi_registers.new_sky\[1\] _02361_
+ vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__mux2_1
X_11707_ clknet_leaf_29_i_clk vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__buf_1
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15475_ _08157_ _08158_ vssd1 vssd1 vccd1 vccd1 _08160_ sky130_fd_sc_hd__and2_1
XFILLER_129_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12687_ _05270_ _05418_ _05419_ _05333_ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__a31o_1
X_17214_ rbzero.wall_tracer.trackDistY\[-7\] _01523_ _01552_ _08539_ vssd1 vssd1 vccd1
+ vccd1 _00564_ sky130_fd_sc_hd__o22a_1
XFILLER_187_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14426_ _04831_ _07111_ _07112_ _07113_ _03490_ vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__a221o_2
X_11638_ rbzero.tex_b1\[57\] rbzero.tex_b1\[56\] _04376_ vssd1 vssd1 vccd1 vccd1 _04419_
+ sky130_fd_sc_hd__mux2_1
X_18194_ rbzero.spi_registers.new_leak\[3\] _02310_ _02316_ _02314_ vssd1 vssd1 vccd1
+ vccd1 _00780_ sky130_fd_sc_hd__o211a_1
XFILLER_200_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17145_ _09231_ _09039_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__or2_1
XFILLER_129_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14357_ _06850_ _05113_ _07044_ _04830_ vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__a211o_1
XFILLER_200_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11569_ rbzero.tex_b0\[19\] rbzero.tex_b0\[18\] _03732_ vssd1 vssd1 vccd1 vccd1 _04351_
+ sky130_fd_sc_hd__mux2_1
XFILLER_144_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13308_ _06058_ _06064_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__xor2_1
X_17076_ _09673_ _09680_ vssd1 vssd1 vccd1 vccd1 _09681_ sky130_fd_sc_hd__and2b_1
Xclkbuf_1_1__f__02734_ clknet_0__02734_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02734_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18956__138 clknet_1_0__leaf__02727_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__inv_2
X_14288_ _06852_ _06679_ _06975_ vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__o21ai_1
XFILLER_170_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16027_ _08359_ _08639_ _08640_ vssd1 vssd1 vccd1 vccd1 _08641_ sky130_fd_sc_hd__a21bo_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13239_ _05472_ _05995_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__nor2_1
XFILLER_170_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17978_ rbzero.pov.spi_buffer\[42\] rbzero.pov.ready_buffer\[42\] _02186_ vssd1 vssd1
+ vccd1 vccd1 _02190_ sky130_fd_sc_hd__mux2_1
X_16929_ _09283_ _09534_ vssd1 vssd1 vccd1 vccd1 _09535_ sky130_fd_sc_hd__xor2_1
XFILLER_133_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19717_ clknet_leaf_3_i_clk _00648_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19648_ clknet_leaf_46_i_clk _00579_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19579_ clknet_leaf_41_i_clk _00510_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20423_ net483 _01354_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20354_ net414 _01285_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20285_ net345 _01216_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10940_ _03666_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__buf_4
XFILLER_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__02754_ clknet_0__02754_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02754_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10871_ _03654_ _03655_ _03656_ vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__mux2_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _05329_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__clkbuf_4
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _06296_ _06344_ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__nor2_1
XFILLER_71_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12541_ _05244_ _05276_ _05297_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__and3_1
XFILLER_185_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_3_0_i_clk clknet_1_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_101_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15260_ _07944_ _07945_ vssd1 vssd1 vccd1 vccd1 _07946_ sky130_fd_sc_hd__nand2_1
XFILLER_8_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12472_ _05087_ _05089_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__nand2_2
XFILLER_185_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19157__319 clknet_1_0__leaf__02747_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__inv_2
XFILLER_71_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14211_ _04838_ rbzero.wall_tracer.stepDistX\[-4\] _06894_ _06898_ vssd1 vssd1 vccd1
+ vccd1 _06899_ sky130_fd_sc_hd__a2bb2o_2
X_11423_ rbzero.tex_g0\[33\] rbzero.tex_g0\[32\] _03699_ vssd1 vssd1 vccd1 vccd1 _04207_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15191_ _07138_ vssd1 vssd1 vccd1 vccd1 _07878_ sky130_fd_sc_hd__clkbuf_4
XFILLER_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_9 _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11354_ rbzero.debug_overlay.playerY\[-8\] _04090_ _04085_ rbzero.debug_overlay.playerY\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__a22o_1
X_14142_ rbzero.wall_tracer.stepDistX\[8\] _06777_ _04833_ vssd1 vssd1 vccd1 vccd1
+ _06836_ sky130_fd_sc_hd__mux2_1
X_10305_ rbzero.tex_b1\[47\] rbzero.tex_b1\[48\] _03210_ vssd1 vssd1 vccd1 vccd1 _03215_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11285_ _04035_ _04049_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__or2_2
X_14073_ rbzero.wall_tracer.visualWallDist\[-3\] _06796_ _06791_ rbzero.wall_tracer.trackDistX\[-3\]
+ _06797_ vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__o221a_1
XFILLER_106_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10236_ rbzero.tex_g0\[17\] rbzero.tex_g0\[16\] _03177_ vssd1 vssd1 vccd1 vccd1 _03179_
+ sky130_fd_sc_hd__mux2_1
X_17901_ _02149_ vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__clkbuf_1
X_13024_ _05494_ _05538_ _05737_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__and3_1
X_18881_ _02708_ vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17832_ _02094_ _02081_ _02085_ vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10167_ rbzero.tex_g0\[49\] rbzero.tex_g0\[48\] _03132_ vssd1 vssd1 vccd1 vccd1 _03142_
+ sky130_fd_sc_hd__mux2_1
XFILLER_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17763_ _02029_ _02027_ _02028_ _03339_ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__o31a_1
X_10098_ _03072_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__clkbuf_4
X_14975_ _06866_ _07661_ _07662_ _06873_ vssd1 vssd1 vccd1 vccd1 _07663_ sky130_fd_sc_hd__o22ai_1
XFILLER_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16714_ _09240_ _09241_ _09321_ vssd1 vssd1 vccd1 vccd1 _09322_ sky130_fd_sc_hd__o21ai_1
X_19502_ clknet_leaf_40_i_clk _00448_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[9\]
+ sky130_fd_sc_hd__dfxtp_4
X_13926_ _06672_ _06674_ _06678_ _05476_ _06629_ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__a221o_2
X_17694_ rbzero.debug_overlay.vplaneX\[-9\] vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__inv_2
XFILLER_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19433_ gpout1.clk_div\[0\] net61 vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__nor2_1
X_16645_ _09016_ _08260_ _09035_ _09014_ vssd1 vssd1 vccd1 vccd1 _09254_ sky130_fd_sc_hd__o22ai_1
XFILLER_35_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13857_ _06560_ _06434_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__xnor2_2
XFILLER_23_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19364_ rbzero.traced_texa\[6\] rbzero.texV\[6\] vssd1 vssd1 vccd1 vccd1 _02844_
+ sky130_fd_sc_hd__or2_1
X_12808_ _05562_ _05563_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__nor2_1
XFILLER_50_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16576_ _09097_ _09185_ vssd1 vssd1 vccd1 vccd1 _09186_ sky130_fd_sc_hd__xnor2_1
X_13788_ _06533_ _06544_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__and2_1
XFILLER_37_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18315_ rbzero.spi_registers.new_other\[3\] rbzero.spi_registers.spi_buffer\[3\]
+ _02388_ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__mux2_1
X_15527_ _08203_ _08210_ vssd1 vssd1 vccd1 vccd1 _08211_ sky130_fd_sc_hd__and2b_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12739_ _05494_ _05488_ _05489_ _05495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__o31a_2
XFILLER_31_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19295_ rbzero.traced_texa\[-5\] rbzero.texV\[-5\] vssd1 vssd1 vccd1 vccd1 _02786_
+ sky130_fd_sc_hd__and2_1
XFILLER_176_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18246_ rbzero.spi_registers.vshift\[2\] _02349_ vssd1 vssd1 vccd1 vccd1 _02352_
+ sky130_fd_sc_hd__or2_1
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15458_ _08020_ _08142_ vssd1 vssd1 vccd1 vccd1 _08143_ sky130_fd_sc_hd__or2_1
XFILLER_124_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19023__198 clknet_1_1__leaf__02734_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__inv_2
X_19097__266 clknet_1_1__leaf__02740_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__inv_2
XFILLER_191_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14409_ _06900_ vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__clkbuf_4
X_18177_ rbzero.spi_registers.new_mapd\[2\] _02289_ _02306_ _02301_ vssd1 vssd1 vccd1
+ vccd1 _00773_ sky130_fd_sc_hd__o211a_1
XFILLER_117_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15389_ _08072_ _08073_ vssd1 vssd1 vccd1 vccd1 _08074_ sky130_fd_sc_hd__nor2_1
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17128_ _01467_ _01471_ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__xnor2_2
XFILLER_190_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09950_ _02983_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__clkbuf_4
X_17059_ _09661_ _09662_ _09663_ vssd1 vssd1 vccd1 vccd1 _09664_ sky130_fd_sc_hd__o21ba_1
XFILLER_131_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__02748_ _02748_ vssd1 vssd1 vccd1 vccd1 clknet_0__02748_ sky130_fd_sc_hd__clkbuf_16
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20070_ clknet_leaf_83_i_clk _01001_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
X_09881_ rbzero.tex_r0\[57\] rbzero.tex_r0\[56\] _02984_ vssd1 vssd1 vccd1 vccd1 _02992_
+ sky130_fd_sc_hd__mux2_1
XFILLER_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20406_ net466 _01337_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20337_ net397 _01268_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 o_gpout[3] sky130_fd_sc_hd__clkbuf_1
XFILLER_1_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11070_ rbzero.map_overlay.i_mapdy\[5\] _03855_ _03840_ vssd1 vssd1 vccd1 vccd1 _03856_
+ sky130_fd_sc_hd__o21a_1
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 o_tex_csb sky130_fd_sc_hd__buf_2
X_20268_ net328 _01199_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10021_ _03065_ vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20199_ net259 _01130_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ _07385_ _07387_ vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__xnor2_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11972_ net2 _04731_ _04725_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__and3_1
XFILLER_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13711_ _06446_ _06466_ _06467_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__a21boi_1
X_10923_ _03662_ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__buf_4
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14691_ _06900_ _06917_ _06939_ _06893_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__o22ai_1
XFILLER_186_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02737_ clknet_0__02737_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02737_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_72_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16430_ _09038_ _09040_ vssd1 vssd1 vccd1 vccd1 _09041_ sky130_fd_sc_hd__xor2_1
XFILLER_32_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13642_ _06231_ _06396_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__xor2_1
X_10854_ rbzero.row_render.texu\[3\] rbzero.row_render.texu\[2\] rbzero.row_render.texu\[1\]
+ _03624_ _03639_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__o32a_1
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _08970_ _08971_ vssd1 vssd1 vccd1 vccd1 _08972_ sky130_fd_sc_hd__nor2_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13573_ _06286_ _06329_ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__nor2_1
XFILLER_169_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10785_ rbzero.traced_texVinit\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _03571_
+ sky130_fd_sc_hd__or2_1
XFILLER_40_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18100_ rbzero.spi_registers.sclk_buffer\[1\] rbzero.spi_registers.sclk_buffer\[0\]
+ _04834_ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__mux2_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15312_ _07880_ _07997_ vssd1 vssd1 vccd1 vccd1 _07998_ sky130_fd_sc_hd__and2_1
XFILLER_12_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12524_ _05220_ _05193_ _05279_ _05259_ _05280_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__o41a_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16292_ _08891_ _08903_ vssd1 vssd1 vccd1 vccd1 _08904_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18031_ _02217_ vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__clkbuf_1
X_15243_ rbzero.debug_overlay.playerY\[-5\] rbzero.debug_overlay.playerX\[-5\] _06851_
+ vssd1 vssd1 vccd1 vccd1 _07930_ sky130_fd_sc_hd__mux2_1
X_12455_ _05126_ _05211_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__xnor2_4
XFILLER_172_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11406_ rbzero.tex_g0\[55\] rbzero.tex_g0\[54\] _04189_ vssd1 vssd1 vccd1 vccd1 _04190_
+ sky130_fd_sc_hd__mux2_1
XFILLER_193_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15174_ _07078_ _06900_ _07039_ _07273_ vssd1 vssd1 vccd1 vccd1 _07861_ sky130_fd_sc_hd__or4_1
XFILLER_165_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12386_ _05141_ _05142_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__xnor2_4
XFILLER_125_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14125_ _06827_ vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11337_ rbzero.debug_overlay.facingX\[10\] _04078_ _04119_ _04121_ vssd1 vssd1 vccd1
+ vccd1 _04122_ sky130_fd_sc_hd__a211o_1
XFILLER_180_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19982_ net211 _00913_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14056_ rbzero.wall_tracer.visualWallDist\[-10\] _03496_ _06785_ rbzero.wall_tracer.trackDistY\[-10\]
+ _03485_ vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__o221a_1
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11268_ gpout0.hpos\[3\] gpout0.hpos\[4\] _04033_ vssd1 vssd1 vccd1 vccd1 _04053_
+ sky130_fd_sc_hd__and3_1
X_13007_ _05761_ _05763_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__xnor2_1
X_10219_ rbzero.tex_g0\[25\] rbzero.tex_g0\[24\] _03166_ vssd1 vssd1 vccd1 vccd1 _03170_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__02433_ clknet_0__02433_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02433_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11199_ rbzero.tex_r1\[24\] _03661_ _03936_ _03983_ vssd1 vssd1 vccd1 vccd1 _03984_
+ sky130_fd_sc_hd__a31o_1
X_19211__368 clknet_1_0__leaf__02752_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__inv_2
X_18864_ _04500_ _04499_ _04508_ _04507_ vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__or4bb_1
X_17815_ _02062_ _02067_ _02077_ _03340_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__a31o_1
X_18795_ rbzero.pov.ready_buffer\[25\] _02644_ _02657_ _02651_ vssd1 vssd1 vccd1 vccd1
+ _01040_ sky130_fd_sc_hd__a211o_1
XFILLER_67_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17746_ _02012_ _02013_ _02010_ _02011_ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__o211ai_1
X_14958_ _07101_ vssd1 vssd1 vccd1 vccd1 _07646_ sky130_fd_sc_hd__buf_2
XFILLER_78_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13909_ _05395_ _06635_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__and2_1
XFILLER_165_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17677_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.wall_tracer.rayAddendX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__nor2_1
X_14889_ _07101_ _07048_ vssd1 vssd1 vccd1 vccd1 _07577_ sky130_fd_sc_hd__nor2_1
X_16628_ _09228_ _09236_ vssd1 vssd1 vccd1 vccd1 _09237_ sky130_fd_sc_hd__and2_1
X_19416_ _01704_ _01709_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__and2b_1
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16559_ _08805_ _09165_ _09168_ vssd1 vssd1 vccd1 vccd1 _09169_ sky130_fd_sc_hd__a21oi_1
X_19347_ _02823_ _02826_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__nand2_1
X_19105__273 clknet_1_0__leaf__02741_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__inv_2
XFILLER_148_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19278_ rbzero.traced_texa\[-8\] rbzero.texV\[-8\] vssd1 vssd1 vccd1 vccd1 _02772_
+ sky130_fd_sc_hd__or2_1
XFILLER_175_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18229_ _02334_ _02340_ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__and2_1
XFILLER_191_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20122_ clknet_leaf_76_i_clk _01053_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
X_09933_ _03019_ vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20053_ clknet_leaf_86_i_clk _00984_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _02981_ _02899_ _02905_ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__or3b_2
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09795_ _02945_ vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10570_ rbzero.debug_overlay.playerX\[1\] _03362_ _03346_ rbzero.debug_overlay.playerY\[2\]
+ _03365_ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__a221o_1
XFILLER_158_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12240_ _04954_ rbzero.wall_tracer.trackDistX\[9\] _04956_ rbzero.wall_tracer.trackDistX\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__o22a_1
XFILLER_147_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12171_ _03375_ _04929_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__nor2_1
XFILLER_135_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11122_ _03849_ _03907_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__nor2_1
XFILLER_150_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11053_ rbzero.debug_overlay.playerX\[3\] vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__inv_2
X_15930_ _08547_ _08548_ _08549_ vssd1 vssd1 vccd1 vccd1 _08550_ sky130_fd_sc_hd__a21oi_1
XFILLER_27_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10004_ _03056_ vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15861_ rbzero.wall_tracer.mapX\[7\] _07825_ vssd1 vssd1 vccd1 vccd1 _08490_ sky130_fd_sc_hd__xor2_1
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ _01882_ _01884_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_0_i_clk i_clk vssd1 vssd1 vccd1 vccd1 clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_77_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14812_ _07456_ _07457_ vssd1 vssd1 vccd1 vccd1 _07500_ sky130_fd_sc_hd__or2_1
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18580_ rbzero.pov.spi_buffer\[58\] rbzero.pov.spi_buffer\[59\] _02499_ vssd1 vssd1
+ vccd1 vccd1 _02509_ sky130_fd_sc_hd__mux2_1
XFILLER_188_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15792_ rbzero.row_render.size\[6\] _08456_ _06717_ _08455_ vssd1 vssd1 vccd1 vccd1
+ _00498_ sky130_fd_sc_hd__a22o_1
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17531_ _01808_ _01811_ _01820_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a21o_1
Xtop_ew_algofoogle_103 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_103/HI zeros[12]
+ sky130_fd_sc_hd__conb_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14743_ _06893_ _06916_ _06939_ _06954_ vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__or4_1
Xtop_ew_algofoogle_114 vssd1 vssd1 vccd1 vccd1 ones[7] top_ew_algofoogle_114/LO sky130_fd_sc_hd__conb_1
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ _04727_ _04728_ net30 vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__mux2_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ rbzero.tex_r0\[23\] rbzero.tex_r0\[22\] _03649_ vssd1 vssd1 vccd1 vccd1 _03692_
+ sky130_fd_sc_hd__mux2_1
X_17462_ _01746_ _01749_ _01747_ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__a21bo_1
XFILLER_83_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14674_ _07359_ _07360_ _07361_ vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__a21oi_1
X_11886_ _04635_ _04659_ _04661_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__a21o_1
XFILLER_17_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16413_ _09020_ _09022_ vssd1 vssd1 vccd1 vccd1 _09024_ sky130_fd_sc_hd__and2_1
X_13625_ _06354_ _06381_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__xnor2_1
X_10837_ _03595_ _03603_ _03622_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__or3_1
X_17393_ rbzero.debug_overlay.playerX\[4\] _01693_ rbzero.wall_tracer.state\[1\] vssd1
+ vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__mux2_1
XFILLER_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19132_ clknet_1_1__leaf__02743_ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__buf_1
XFILLER_201_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16344_ _08831_ _08721_ vssd1 vssd1 vccd1 vccd1 _08956_ sky130_fd_sc_hd__or2b_1
XFILLER_185_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13556_ _06173_ _06262_ _06261_ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__nand3_1
XFILLER_73_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10768_ rbzero.traced_texVinit\[2\] rbzero.texV\[2\] rbzero.texV\[1\] rbzero.traced_texVinit\[1\]
+ _03553_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__a221o_1
XFILLER_200_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12507_ _05197_ _05257_ _05254_ _05263_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__or4_1
Xclkbuf_1_0_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_1_0_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_16275_ _08768_ _08885_ _08886_ vssd1 vssd1 vccd1 vccd1 _08887_ sky130_fd_sc_hd__o21ai_1
XFILLER_160_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13487_ _06241_ _06243_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10699_ _03488_ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__clkbuf_4
X_18014_ rbzero.pov.spi_buffer\[59\] rbzero.pov.ready_buffer\[59\] _02208_ vssd1 vssd1
+ vccd1 vccd1 _02209_ sky130_fd_sc_hd__mux2_1
XFILLER_195_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15226_ _07910_ _07912_ vssd1 vssd1 vccd1 vccd1 _07913_ sky130_fd_sc_hd__xor2_1
XFILLER_145_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12438_ _05133_ _05147_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__nor2_1
XFILLER_154_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15157_ _07842_ _07843_ vssd1 vssd1 vccd1 vccd1 _07844_ sky130_fd_sc_hd__or2_1
X_12369_ _05124_ _05125_ _05072_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__mux2_2
XFILLER_114_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14108_ _06818_ vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19965_ net194 _00896_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[45\] sky130_fd_sc_hd__dfxtp_1
X_15088_ _07727_ _07775_ vssd1 vssd1 vccd1 vccd1 _07776_ sky130_fd_sc_hd__xnor2_1
X_19135__299 clknet_1_0__leaf__02745_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__inv_2
XFILLER_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14039_ _06774_ _06776_ vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__nand2_1
XFILLER_141_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19896_ clknet_leaf_19_i_clk _00827_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18847_ rbzero.debug_overlay.vplaneY\[-4\] _02634_ vssd1 vssd1 vccd1 vccd1 _02686_
+ sky130_fd_sc_hd__and2_1
XFILLER_67_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18778_ rbzero.pov.ready_buffer\[39\] _02644_ _02648_ _02559_ vssd1 vssd1 vccd1 vccd1
+ _01032_ sky130_fd_sc_hd__a211o_1
XFILLER_36_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17729_ _08458_ _01989_ _01990_ _01999_ vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__a31o_1
XFILLER_36_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20105_ clknet_leaf_88_i_clk _01036_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[10\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_3_2_0_i_clk clknet_2_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09916_ _03010_ vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20036_ clknet_leaf_0_i_clk _00967_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09847_ _02972_ vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__clkbuf_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09778_ _02936_ vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__clkbuf_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11740_ gpout0.clk_div\[1\] _04515_ _04513_ _04517_ vssd1 vssd1 vccd1 vccd1 _04518_
+ sky130_fd_sc_hd__a31o_2
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11671_ rbzero.tex_b1\[11\] rbzero.tex_b1\[10\] _04376_ vssd1 vssd1 vccd1 vccd1 _04452_
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ _05549_ _06055_ _05610_ _06061_ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_168_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10622_ _03415_ _03416_ _03417_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__or3_1
X_14390_ _06908_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0__f__02436_ clknet_0__02436_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02436_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_139_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13341_ _06097_ _06055_ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__nor2_2
XFILLER_195_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10553_ _03342_ _03343_ rbzero.map_rom.i_row\[4\] _03344_ _03348_ vssd1 vssd1 vccd1
+ vccd1 _03349_ sky130_fd_sc_hd__a221o_1
XFILLER_154_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16060_ _07661_ _08018_ _08392_ vssd1 vssd1 vccd1 vccd1 _08674_ sky130_fd_sc_hd__o21ai_1
XFILLER_127_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13272_ _05972_ _06005_ _06028_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__o21ai_1
XFILLER_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10484_ _03308_ vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15011_ _07479_ _07573_ _07696_ _07698_ vssd1 vssd1 vccd1 vccd1 _07699_ sky130_fd_sc_hd__a22o_2
XFILLER_170_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12223_ rbzero.wall_tracer.trackDistY\[-2\] vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__inv_2
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12154_ _04911_ _04915_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__nand2_1
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11105_ gpout0.vpos\[2\] rbzero.debug_overlay.playerY\[-1\] vssd1 vssd1 vccd1 vccd1
+ _03891_ sky130_fd_sc_hd__xnor2_1
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19750_ clknet_leaf_92_i_clk _00681_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16962_ _09433_ _09566_ _09567_ vssd1 vssd1 vccd1 vccd1 _09568_ sky130_fd_sc_hd__o21ai_1
X_12085_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] vssd1
+ vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__or2_1
XFILLER_150_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18701_ _02588_ _02590_ _02591_ _02319_ vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__a211oi_1
X_11036_ _03726_ _03768_ _03769_ _03821_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__o31a_1
X_15913_ _08526_ _08527_ _08528_ vssd1 vssd1 vccd1 vccd1 _08535_ sky130_fd_sc_hd__o21bai_1
X_16893_ _09476_ _09499_ vssd1 vssd1 vccd1 vccd1 _09500_ sky130_fd_sc_hd__xnor2_1
X_19681_ clknet_leaf_80_i_clk _00612_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18632_ _02261_ _02411_ vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__and2_1
X_15844_ _03362_ _07936_ _08473_ vssd1 vssd1 vccd1 vccd1 _08474_ sky130_fd_sc_hd__o21ai_1
XFILLER_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15775_ _03508_ vssd1 vssd1 vccd1 vccd1 _08447_ sky130_fd_sc_hd__buf_4
X_18563_ _02500_ vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__clkbuf_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _05707_ _05734_ _05739_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__and3_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _07066_ _07413_ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__xnor2_1
X_17514_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.debug_overlay.vplaneY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__or2_1
XFILLER_45_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18494_ rbzero.pov.spi_buffer\[17\] rbzero.pov.spi_buffer\[18\] _02455_ vssd1 vssd1
+ vccd1 vccd1 _02464_ sky130_fd_sc_hd__mux2_1
X_11938_ net39 _04665_ _04669_ net49 vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__a22o_1
XFILLER_33_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17445_ _01739_ _01740_ _03486_ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__a21oi_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14657_ _06908_ _07147_ vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__or2_1
X_11869_ net10 net11 net12 vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__a21o_1
XFILLER_20_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13608_ _06316_ _06315_ _06173_ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__a21o_1
XFILLER_60_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17376_ _03395_ _01680_ _08507_ vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__mux2_1
X_14588_ _07275_ vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__inv_2
XFILLER_159_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16327_ _08812_ _08813_ _08815_ vssd1 vssd1 vccd1 vccd1 _08939_ sky130_fd_sc_hd__o21a_1
XFILLER_173_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13539_ _05503_ _06071_ vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__nor2_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16258_ _08868_ _08869_ vssd1 vssd1 vccd1 vccd1 _08870_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15209_ _03492_ rbzero.wall_tracer.stepDistY\[6\] _04949_ vssd1 vssd1 vccd1 vccd1
+ _07896_ sky130_fd_sc_hd__a21o_1
XFILLER_173_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16189_ _08798_ _08801_ vssd1 vssd1 vccd1 vccd1 _08802_ sky130_fd_sc_hd__xnor2_1
X_19217__374 clknet_1_1__leaf__02752_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__inv_2
XFILLER_99_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19948_ net177 _00879_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19879_ clknet_leaf_21_i_clk _00810_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_63_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_78_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20019_ clknet_leaf_94_i_clk _00950_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12910_ _05493_ _05536_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__nor2_1
XFILLER_98_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13890_ _06588_ _05395_ _06609_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__and3_1
XFILLER_101_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12841_ _05588_ _05597_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__xnor2_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_16_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _08131_ _08135_ _08132_ vssd1 vssd1 vccd1 vccd1 _08244_ sky130_fd_sc_hd__a21bo_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12772_ _05525_ _05518_ _05528_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__or3b_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _07178_ vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__clkbuf_4
XFILLER_14_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _03906_ _04499_ _03909_ _04500_ _04494_ _04487_ vssd1 vssd1 vccd1 vccd1 _04501_
+ sky130_fd_sc_hd__mux4_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _08174_ _08175_ vssd1 vssd1 vccd1 vccd1 _08176_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ rbzero.wall_tracer.trackDistY\[-4\] rbzero.wall_tracer.stepDistY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__or2_1
XFILLER_14_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _06733_ _07103_ _06738_ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__a21o_1
XFILLER_175_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11654_ rbzero.tex_b1\[31\] rbzero.tex_b1\[30\] _04376_ vssd1 vssd1 vccd1 vccd1 _04435_
+ sky130_fd_sc_hd__mux2_1
XFILLER_168_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17161_ _01495_ _01504_ vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10605_ _03373_ _03352_ _03399_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__o21ai_1
XFILLER_196_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14373_ _07054_ _07059_ vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__nand2_1
XFILLER_11_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11585_ rbzero.tex_b0\[11\] _04155_ _04156_ _03659_ vssd1 vssd1 vccd1 vccd1 _04367_
+ sky130_fd_sc_hd__a31o_1
XFILLER_11_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16112_ _08633_ _08722_ _08724_ vssd1 vssd1 vccd1 vccd1 _08725_ sky130_fd_sc_hd__a21oi_4
XFILLER_156_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13324_ _05962_ _06056_ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__and2_1
XFILLER_70_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17092_ _09595_ _09694_ _09695_ vssd1 vssd1 vccd1 vccd1 _09697_ sky130_fd_sc_hd__or3b_1
XFILLER_183_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__02750_ clknet_0__02750_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02750_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_156_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10536_ _03335_ vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16043_ _08638_ _08386_ _08656_ vssd1 vssd1 vccd1 vccd1 _08657_ sky130_fd_sc_hd__a21o_1
X_13255_ _05953_ _06007_ _06010_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__nor3_1
X_10467_ _03299_ vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12206_ _04964_ rbzero.wall_tracer.trackDistX\[-1\] _04967_ vssd1 vssd1 vccd1 vccd1
+ _04968_ sky130_fd_sc_hd__o21ai_1
X_13186_ _05888_ _05908_ _05941_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__and3_1
X_10398_ _03263_ vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19802_ clknet_leaf_15_i_clk _00733_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12137_ _04857_ _04864_ _04852_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__nand3_1
X_17994_ _02198_ vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19733_ clknet_leaf_93_i_clk _00664_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16945_ _09549_ _09550_ vssd1 vssd1 vccd1 vccd1 _09551_ sky130_fd_sc_hd__and2_1
X_12068_ _04835_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11019_ rbzero.row_render.size\[3\] _03772_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__nand2_1
X_19664_ clknet_leaf_4_i_clk _00595_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_16876_ _09142_ _08889_ vssd1 vssd1 vccd1 vccd1 _09483_ sky130_fd_sc_hd__nor2_1
XFILLER_77_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18615_ net51 rbzero.pov.ss_buffer\[0\] _03337_ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__mux2_1
XFILLER_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827_ rbzero.traced_texa\[6\] _08463_ _08462_ rbzero.wall_tracer.visualWallDist\[6\]
+ vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__a22o_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19595_ clknet_leaf_44_i_clk _00526_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18546_ _02491_ vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__clkbuf_1
X_15758_ _02981_ _03506_ vssd1 vssd1 vccd1 vccd1 _08439_ sky130_fd_sc_hd__nor2_8
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14709_ _06949_ _06977_ _07005_ _06966_ vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__o22a_1
X_15689_ _08370_ _08371_ vssd1 vssd1 vccd1 vccd1 _08372_ sky130_fd_sc_hd__xor2_1
X_18477_ _02443_ vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__clkbuf_4
XFILLER_127_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17428_ rbzero.wall_tracer.rayAddendY\[-4\] _00013_ _01721_ _01725_ vssd1 vssd1 vccd1
+ vccd1 _00605_ sky130_fd_sc_hd__o22a_1
XFILLER_193_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17359_ rbzero.spi_registers.new_mapd\[8\] rbzero.spi_registers.spi_buffer\[8\] _01663_
+ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__mux2_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20370_ net430 _01301_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18933__117 clknet_1_0__leaf__02725_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__inv_2
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11370_ rbzero.tex_g0\[17\] rbzero.tex_g0\[16\] _03663_ vssd1 vssd1 vccd1 vccd1 _04154_
+ sky130_fd_sc_hd__mux2_1
XFILLER_180_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10321_ _03223_ vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20499_ clknet_leaf_41_i_clk _01430_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_152_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13040_ _05791_ _05795_ _05796_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__o21ai_1
X_10252_ rbzero.tex_g0\[9\] rbzero.tex_g0\[8\] _03177_ vssd1 vssd1 vccd1 vccd1 _03187_
+ sky130_fd_sc_hd__mux2_1
XFILLER_140_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10183_ rbzero.tex_g0\[42\] rbzero.tex_g0\[41\] _03144_ vssd1 vssd1 vccd1 vccd1 _03151_
+ sky130_fd_sc_hd__mux2_1
XFILLER_132_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14991_ _07265_ _07213_ vssd1 vssd1 vccd1 vccd1 _07679_ sky130_fd_sc_hd__nand2_1
XFILLER_87_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16730_ _07766_ _09231_ _09229_ _08899_ vssd1 vssd1 vccd1 vccd1 _09338_ sky130_fd_sc_hd__o22ai_1
X_13942_ _05447_ _06610_ _06692_ _06675_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__a22o_1
XFILLER_120_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16661_ _08245_ _08678_ vssd1 vssd1 vccd1 vccd1 _09270_ sky130_fd_sc_hd__nor2_1
XFILLER_35_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13873_ _06629_ vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__clkbuf_4
XFILLER_35_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15612_ _08294_ _08295_ vssd1 vssd1 vccd1 vccd1 _08296_ sky130_fd_sc_hd__and2_1
XFILLER_62_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12824_ _05577_ _05579_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__nand2_1
XFILLER_74_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19380_ _02854_ _02855_ _02856_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__nand3_1
X_16592_ _09200_ _09201_ vssd1 vssd1 vccd1 vccd1 _09202_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15543_ _07984_ _07857_ vssd1 vssd1 vccd1 vccd1 _08227_ sky130_fd_sc_hd__nor2_1
X_18331_ _02107_ _01658_ _02907_ _02399_ vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__and4b_1
X_12755_ _05510_ _05511_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__and2b_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _03471_ _04475_ _04485_ net69 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__o22ai_4
X_18262_ _02362_ vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__clkbuf_1
XFILLER_148_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15474_ _08157_ _08158_ vssd1 vssd1 vccd1 vccd1 _08159_ sky130_fd_sc_hd__nor2_1
XFILLER_188_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _05310_ _05323_ _05434_ _05439_ _05442_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__a32oi_4
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14425_ _06850_ _05143_ _04830_ vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__a21oi_1
X_17213_ _01534_ _01550_ _01551_ _01526_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__a31o_1
X_11637_ _04416_ _04417_ _03656_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__mux2_1
XFILLER_128_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18193_ rbzero.floor_leak\[3\] _02311_ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__or2_1
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17144_ _01482_ _01487_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14356_ _06849_ _04896_ vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__nor2_1
X_11568_ rbzero.tex_b0\[17\] rbzero.tex_b0\[16\] _04189_ vssd1 vssd1 vccd1 vccd1 _04350_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13307_ _06059_ _06063_ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__xnor2_1
X_17075_ _09674_ _09679_ vssd1 vssd1 vccd1 vccd1 _09680_ sky130_fd_sc_hd__xor2_1
Xclkbuf_1_1__f__02733_ clknet_0__02733_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02733_
+ sky130_fd_sc_hd__clkbuf_16
X_10519_ rbzero.tex_b0\[10\] rbzero.tex_b0\[9\] _03324_ vssd1 vssd1 vccd1 vccd1 _03327_
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14287_ _04830_ _06974_ _06859_ vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__o21a_1
X_11499_ rbzero.tex_g1\[63\] _03729_ _03730_ _03661_ vssd1 vssd1 vccd1 vccd1 _04282_
+ sky130_fd_sc_hd__a31o_1
XFILLER_143_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16026_ _06856_ _06874_ _07141_ _07092_ vssd1 vssd1 vccd1 vccd1 _08640_ sky130_fd_sc_hd__or4_2
X_13238_ _05994_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__clkbuf_4
XFILLER_112_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13169_ _05433_ _05517_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__or2_1
XFILLER_151_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17977_ _02189_ vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19716_ clknet_leaf_3_i_clk _00647_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16928_ _09470_ _09533_ vssd1 vssd1 vccd1 vccd1 _09534_ sky130_fd_sc_hd__xor2_2
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19647_ clknet_leaf_45_i_clk _00578_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19028__203 clknet_1_0__leaf__02734_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__inv_2
X_16859_ _07992_ _08803_ vssd1 vssd1 vccd1 vccd1 _09466_ sky130_fd_sc_hd__nor2_1
XFILLER_92_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18442__81 clknet_1_0__leaf__02439_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__inv_2
XFILLER_129_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19578_ clknet_leaf_37_i_clk _00509_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
X_18529_ _02482_ vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20422_ net482 _01353_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20353_ net413 _01284_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19074__245 clknet_1_1__leaf__02738_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__inv_2
XFILLER_175_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20284_ net344 _01215_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__02753_ clknet_0__02753_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02753_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_83_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10870_ _03635_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__buf_6
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12540_ _05286_ _05290_ _05293_ _05296_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__nor4b_4
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12471_ _05094_ _05227_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__xor2_2
XFILLER_200_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14210_ _06852_ _06705_ _06897_ vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__o21ai_1
XFILLER_184_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11422_ _04198_ _04201_ _04205_ _03721_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__a211o_1
X_15190_ _07100_ vssd1 vssd1 vccd1 vccd1 _07877_ sky130_fd_sc_hd__clkbuf_4
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14141_ _06835_ vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__clkbuf_1
X_11353_ rbzero.debug_overlay.playerY\[1\] _04066_ _04068_ rbzero.debug_overlay.playerY\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__a22o_1
XFILLER_192_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10304_ _03214_ vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__clkbuf_1
X_14072_ rbzero.wall_tracer.trackDistY\[-4\] _06786_ _06799_ vssd1 vssd1 vccd1 vccd1
+ _00435_ sky130_fd_sc_hd__o21a_1
X_11284_ _04064_ _04066_ _04068_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__or3_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17900_ rbzero.pov.spi_buffer\[5\] rbzero.pov.ready_buffer\[5\] _02143_ vssd1 vssd1
+ vccd1 vccd1 _02149_ sky130_fd_sc_hd__mux2_1
X_13023_ _05494_ _05538_ _05737_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__a21o_1
X_10235_ _03178_ vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__clkbuf_1
X_18880_ _02287_ _02706_ _02707_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__and3b_1
XFILLER_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17831_ _02001_ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__inv_2
X_10166_ _03141_ vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17762_ _02027_ _02028_ _02029_ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__o21ai_1
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10097_ _03105_ vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__clkbuf_1
X_14974_ _07646_ vssd1 vssd1 vccd1 vccd1 _07662_ sky130_fd_sc_hd__buf_2
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19501_ clknet_leaf_46_i_clk _00447_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[8\]
+ sky130_fd_sc_hd__dfxtp_4
X_16713_ _09226_ _09242_ vssd1 vssd1 vccd1 vccd1 _09321_ sky130_fd_sc_hd__or2b_1
XFILLER_48_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13925_ _06675_ _06677_ vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__and2_1
X_17693_ _01961_ _01962_ _01964_ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a21o_1
XFILLER_48_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19432_ _02885_ _02886_ rbzero.wall_tracer.rayAddendX\[-6\] _08449_ vssd1 vssd1 vccd1
+ vccd1 _01448_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16644_ _07494_ _08229_ _08260_ _08018_ vssd1 vssd1 vccd1 vccd1 _09253_ sky130_fd_sc_hd__or4_1
X_13856_ _06610_ _06612_ vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__or2_1
XFILLER_90_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12807_ _05562_ _05563_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__xor2_1
XFILLER_90_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19363_ rbzero.texV\[5\] _02762_ _02709_ _02843_ vssd1 vssd1 vccd1 vccd1 _01422_
+ sky130_fd_sc_hd__a22o_1
X_16575_ _09183_ _09184_ vssd1 vssd1 vccd1 vccd1 _09185_ sky130_fd_sc_hd__and2b_1
X_13787_ _05805_ _06156_ _06532_ vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__o21ai_1
XFILLER_43_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10999_ rbzero.row_render.size\[2\] _03783_ _03499_ rbzero.row_render.size\[1\] _03784_
+ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__o221a_1
XFILLER_16_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18314_ _02391_ vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__clkbuf_1
X_15526_ _08208_ _08209_ vssd1 vssd1 vccd1 vccd1 _08210_ sky130_fd_sc_hd__xnor2_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _05404_ _05425_ _05449_ _05443_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__a211o_4
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19294_ rbzero.traced_texa\[-5\] rbzero.texV\[-5\] vssd1 vssd1 vccd1 vccd1 _02785_
+ sky130_fd_sc_hd__nor2_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18245_ rbzero.spi_registers.new_vshift\[1\] _02348_ _02351_ _02314_ vssd1 vssd1
+ vccd1 vccd1 _00796_ sky130_fd_sc_hd__o211a_1
X_15457_ _07195_ _04949_ _03493_ _08141_ vssd1 vssd1 vccd1 vccd1 _08142_ sky130_fd_sc_hd__or4_2
XFILLER_198_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12669_ _05367_ _05405_ _05407_ _05274_ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__a211o_1
X_14408_ _07080_ _07093_ _07095_ vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__o21a_1
XFILLER_198_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15388_ _07269_ _07961_ _08071_ _07011_ vssd1 vssd1 vccd1 vccd1 _08073_ sky130_fd_sc_hd__o22a_1
XFILLER_129_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18176_ rbzero.mapdxw\[0\] _02291_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__or2_1
XFILLER_190_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17127_ _01468_ _01470_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__xor2_1
X_14339_ rbzero.debug_overlay.playerY\[-2\] _06980_ rbzero.debug_overlay.playerY\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _07027_ sky130_fd_sc_hd__o21ai_1
XFILLER_143_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17058_ _08896_ _07961_ _08071_ _08899_ vssd1 vssd1 vccd1 vccd1 _09663_ sky130_fd_sc_hd__o22a_1
XFILLER_144_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16009_ _08621_ _08622_ vssd1 vssd1 vccd1 vccd1 _08623_ sky130_fd_sc_hd__xor2_1
XFILLER_131_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__02747_ _02747_ vssd1 vssd1 vccd1 vccd1 clknet_0__02747_ sky130_fd_sc_hd__clkbuf_16
XFILLER_83_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09880_ _02991_ vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__clkbuf_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20405_ net465 _01336_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18939__123 clknet_1_0__leaf__02725_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__inv_2
XFILLER_174_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20336_ net396 _01267_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 o_gpout[4] sky130_fd_sc_hd__clkbuf_1
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 o_tex_oeb0 sky130_fd_sc_hd__buf_2
X_20267_ net327 _01198_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10020_ rbzero.tex_g1\[54\] rbzero.tex_g1\[55\] _03061_ vssd1 vssd1 vccd1 vccd1 _03065_
+ sky130_fd_sc_hd__mux2_1
XFILLER_131_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20198_ net258 _01129_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ net51 _04731_ _04732_ _04532_ _04744_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__a221o_1
XFILLER_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13710_ _06447_ _06448_ _06465_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__nand3_1
XFILLER_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10922_ _03706_ _03707_ _03693_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__mux2_1
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14690_ _06917_ _06939_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__nor2_1
XFILLER_186_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18985__165 clknet_1_0__leaf__02729_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__inv_2
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__02736_ clknet_0__02736_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02736_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18421__62 clknet_1_1__leaf__02437_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__inv_2
XFILLER_60_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13641_ _06357_ _06378_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__xnor2_1
X_10853_ _03634_ _03635_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__nand2_1
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _08879_ _08968_ _08969_ vssd1 vssd1 vccd1 vccd1 _08971_ sky130_fd_sc_hd__and3_1
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13572_ _06304_ _06327_ _06328_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__a21oi_1
XFILLER_201_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10784_ _03568_ _03569_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__xnor2_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15311_ _07530_ _07137_ vssd1 vssd1 vccd1 vccd1 _07997_ sky130_fd_sc_hd__nor2_1
XFILLER_13_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12523_ _05189_ _05192_ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__or2_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16291_ _08901_ _08902_ vssd1 vssd1 vccd1 vccd1 _08903_ sky130_fd_sc_hd__nor2_1
XFILLER_185_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18030_ rbzero.pov.spi_buffer\[67\] rbzero.pov.ready_buffer\[67\] _02208_ vssd1 vssd1
+ vccd1 vccd1 _02217_ sky130_fd_sc_hd__mux2_1
X_15242_ _07830_ _07928_ vssd1 vssd1 vccd1 vccd1 _07929_ sky130_fd_sc_hd__xnor2_4
X_12454_ _05120_ _05199_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__nand2_1
XFILLER_173_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11405_ _04188_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__buf_6
X_15173_ _07078_ _07039_ vssd1 vssd1 vccd1 vccd1 _07860_ sky130_fd_sc_hd__or2_1
X_12385_ _05051_ _05054_ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__nand2_2
XFILLER_181_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14124_ rbzero.wall_tracer.stepDistX\[-1\] _06726_ _06825_ vssd1 vssd1 vccd1 vccd1
+ _06827_ sky130_fd_sc_hd__mux2_1
XFILLER_197_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11336_ rbzero.debug_overlay.facingX\[-3\] _04092_ _04056_ rbzero.debug_overlay.facingX\[-2\]
+ _04120_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__a221o_1
XFILLER_193_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19981_ net210 _00912_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18932_ clknet_1_0__leaf__02440_ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__buf_1
X_14055_ rbzero.wall_tracer.trackDistY\[-11\] _06786_ _06789_ vssd1 vssd1 vccd1 vccd1
+ _00428_ sky130_fd_sc_hd__o21a_1
X_11267_ _03504_ _03514_ _04045_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__or3b_2
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13006_ _05722_ _05724_ _05762_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__a21oi_1
X_10218_ _03169_ vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__clkbuf_1
X_18863_ _02258_ _02694_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__nand2_1
X_11198_ rbzero.tex_r1\[25\] _03660_ _03768_ _03670_ vssd1 vssd1 vccd1 vccd1 _03983_
+ sky130_fd_sc_hd__a31o_1
XFILLER_121_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17814_ _02062_ _02067_ _02077_ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__a21oi_1
XFILLER_79_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10149_ rbzero.tex_g0\[58\] rbzero.tex_g0\[57\] _03132_ vssd1 vssd1 vccd1 vccd1 _03133_
+ sky130_fd_sc_hd__mux2_1
X_18794_ rbzero.debug_overlay.facingY\[-6\] _02645_ vssd1 vssd1 vccd1 vccd1 _02657_
+ sky130_fd_sc_hd__and2_1
XFILLER_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17745_ _02010_ _02011_ _02012_ _02013_ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__a211o_1
XFILLER_36_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14957_ _07634_ _07644_ vssd1 vssd1 vccd1 vccd1 _07645_ sky130_fd_sc_hd__nand2_1
XFILLER_63_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13908_ _05421_ _06640_ _06645_ _05372_ _06637_ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__o221a_1
X_17676_ rbzero.wall_tracer.rayAddendX\[-3\] _00013_ _01947_ _01950_ vssd1 vssd1 vccd1
+ vccd1 _00628_ sky130_fd_sc_hd__o22a_1
X_14888_ _07547_ _07566_ vssd1 vssd1 vccd1 vccd1 _07576_ sky130_fd_sc_hd__xor2_1
X_19415_ rbzero.wall_tracer.rayAddendY\[-8\] _02868_ _08454_ _02875_ vssd1 vssd1 vccd1
+ vccd1 _01442_ sky130_fd_sc_hd__a22o_1
X_16627_ _09234_ _09235_ vssd1 vssd1 vccd1 vccd1 _09236_ sky130_fd_sc_hd__xnor2_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13839_ _05696_ _06098_ _06081_ _06097_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__a211o_1
XFILLER_189_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19346_ rbzero.traced_texa\[3\] rbzero.texV\[3\] vssd1 vssd1 vccd1 vccd1 _02829_
+ sky130_fd_sc_hd__nand2_1
X_16558_ _08807_ _09167_ vssd1 vssd1 vccd1 vccd1 _09168_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15509_ _07265_ _08069_ vssd1 vssd1 vccd1 vccd1 _08193_ sky130_fd_sc_hd__nor2_1
XFILLER_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19277_ rbzero.texV\[-9\] _02675_ _02709_ _02771_ vssd1 vssd1 vccd1 vccd1 _01408_
+ sky130_fd_sc_hd__a22o_1
X_16489_ _09029_ _09006_ vssd1 vssd1 vccd1 vccd1 _09099_ sky130_fd_sc_hd__or2b_1
XFILLER_176_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18228_ rbzero.color_floor\[2\] rbzero.spi_registers.new_floor\[2\] _02335_ vssd1
+ vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__mux2_1
XFILLER_191_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18159_ rbzero.map_overlay.i_mapdx\[4\] _02292_ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__or2_1
XFILLER_117_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09932_ rbzero.tex_r0\[33\] rbzero.tex_r0\[32\] _03017_ vssd1 vssd1 vccd1 vccd1 _03019_
+ sky130_fd_sc_hd__mux2_1
XFILLER_144_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20121_ clknet_leaf_77_i_clk _01052_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20052_ clknet_leaf_85_i_clk _00983_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09863_ _02906_ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__clkinv_8
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ rbzero.tex_r1\[32\] rbzero.tex_r1\[33\] _02943_ vssd1 vssd1 vccd1 vccd1 _02945_
+ sky130_fd_sc_hd__mux2_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19186__346 clknet_1_0__leaf__02749_ vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__inv_2
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12170_ rbzero.map_rom.i_row\[4\] _04929_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__xnor2_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11121_ gpout0.vpos\[7\] gpout0.vpos\[6\] vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__nand2_1
XFILLER_162_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20319_ net379 _01250_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_122_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11052_ _03466_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__buf_4
XFILLER_104_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10003_ rbzero.tex_g1\[62\] rbzero.tex_g1\[63\] _02976_ vssd1 vssd1 vccd1 vccd1 _03056_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15860_ _08483_ _08484_ _08488_ _08489_ rbzero.wall_tracer.mapX\[6\] vssd1 vssd1
+ vccd1 vccd1 _00533_ sky130_fd_sc_hd__a32o_1
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14811_ _07446_ _07460_ vssd1 vssd1 vccd1 vccd1 _07499_ sky130_fd_sc_hd__xnor2_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ rbzero.row_render.size\[5\] _08456_ _06712_ _08455_ vssd1 vssd1 vccd1 vccd1
+ _00497_ sky130_fd_sc_hd__a22o_1
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _01818_ _01819_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__nand2_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11954_ gpout0.hpos\[0\] _03527_ _03526_ _04020_ net27 net28 vssd1 vssd1 vccd1 vccd1
+ _04728_ sky130_fd_sc_hd__mux4_1
XFILLER_18_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14742_ _06917_ _06939_ _06969_ _06893_ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__o22a_1
Xtop_ew_algofoogle_104 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_104/HI zeros[13]
+ sky130_fd_sc_hd__conb_1
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_115 vssd1 vssd1 vccd1 vccd1 ones[8] top_ew_algofoogle_115/LO sky130_fd_sc_hd__conb_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ rbzero.tex_r0\[21\] rbzero.tex_r0\[20\] _03690_ vssd1 vssd1 vccd1 vccd1 _03691_
+ sky130_fd_sc_hd__mux2_1
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17461_ _01745_ _01750_ _01751_ _01755_ vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__a31o_1
XFILLER_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14673_ _07341_ _07358_ vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__nor2_1
XFILLER_189_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11885_ _04623_ _04660_ _04647_ net13 vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__a211o_1
XFILLER_83_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16412_ _09020_ _09022_ vssd1 vssd1 vccd1 vccd1 _09023_ sky130_fd_sc_hd__nor2_1
X_13624_ _06355_ _06380_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__xor2_1
X_10836_ _03593_ _03594_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__and2_1
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17392_ _08471_ _08480_ vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__xor2_1
XFILLER_198_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16343_ _08719_ _08720_ _08831_ _08711_ vssd1 vssd1 vccd1 vccd1 _08955_ sky130_fd_sc_hd__a31o_1
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13555_ _06291_ _06311_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10767_ rbzero.traced_texVinit\[1\] rbzero.texV\[1\] rbzero.texV\[0\] rbzero.traced_texVinit\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__o211a_1
XFILLER_158_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12506_ _05220_ _05193_ _05259_ _05262_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__or4_1
XFILLER_201_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16274_ _06858_ _07012_ _07878_ _08252_ vssd1 vssd1 vccd1 vccd1 _08886_ sky130_fd_sc_hd__or4_1
XFILLER_160_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13486_ _06152_ _06242_ vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__and2_1
XFILLER_160_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10698_ _03487_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__clkbuf_4
XFILLER_200_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15225_ _07741_ _07770_ _07911_ vssd1 vssd1 vccd1 vccd1 _07912_ sky130_fd_sc_hd__a21oi_1
X_18013_ _02141_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__buf_4
X_12437_ _05065_ _05069_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__nand2_1
XFILLER_173_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15156_ _07709_ _07834_ _07841_ vssd1 vssd1 vccd1 vccd1 _07843_ sky130_fd_sc_hd__a21oi_1
XFILLER_153_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12368_ rbzero.wall_tracer.visualWallDist\[-7\] _04890_ rbzero.wall_tracer.rcp_sel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__mux2_1
XFILLER_141_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14107_ rbzero.wall_tracer.stepDistX\[-9\] _06658_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _06818_ sky130_fd_sc_hd__mux2_1
XFILLER_181_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11319_ rbzero.debug_overlay.vplaneX\[-3\] _04092_ _04101_ _04103_ vssd1 vssd1 vccd1
+ vccd1 _04104_ sky130_fd_sc_hd__a211o_1
XFILLER_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19964_ net193 _00895_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[44\] sky130_fd_sc_hd__dfxtp_1
X_15087_ _07773_ _07774_ vssd1 vssd1 vccd1 vccd1 _07775_ sky130_fd_sc_hd__and2b_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12299_ rbzero.debug_overlay.facingX\[-1\] rbzero.wall_tracer.rayAddendX\[7\] vssd1
+ vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__and2_1
X_14038_ _05210_ _05278_ _05322_ _06731_ _06775_ vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__a221o_1
XFILLER_113_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19895_ clknet_leaf_19_i_clk _00826_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18846_ rbzero.pov.ready_buffer\[4\] _02666_ _02685_ _02675_ vssd1 vssd1 vccd1 vccd1
+ _01063_ sky130_fd_sc_hd__a211o_1
XFILLER_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18777_ rbzero.debug_overlay.facingX\[-3\] _02645_ vssd1 vssd1 vccd1 vccd1 _02648_
+ sky130_fd_sc_hd__and2_1
X_15989_ _08601_ _08602_ vssd1 vssd1 vccd1 vccd1 _08603_ sky130_fd_sc_hd__nor2_1
XFILLER_82_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17728_ _01722_ _01997_ _01998_ _08448_ rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__a32o_1
XFILLER_24_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17659_ _01916_ _01929_ _01917_ vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__o21ai_1
XFILLER_23_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18400__43 clknet_1_1__leaf__02435_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__inv_2
XFILLER_149_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19329_ _02811_ _02812_ _02806_ _02810_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__a211o_1
XFILLER_176_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20104_ clknet_leaf_89_i_clk _01035_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_09915_ rbzero.tex_r0\[41\] rbzero.tex_r0\[40\] _03006_ vssd1 vssd1 vccd1 vccd1 _03010_
+ sky130_fd_sc_hd__mux2_1
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09846_ rbzero.tex_r1\[7\] rbzero.tex_r1\[8\] _02965_ vssd1 vssd1 vccd1 vccd1 _02972_
+ sky130_fd_sc_hd__mux2_1
X_20035_ clknet_leaf_0_i_clk _00966_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09777_ rbzero.tex_r1\[40\] rbzero.tex_r1\[41\] _02932_ vssd1 vssd1 vccd1 vccd1 _02936_
+ sky130_fd_sc_hd__mux2_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ rbzero.tex_b1\[9\] rbzero.tex_b1\[8\] _04376_ vssd1 vssd1 vccd1 vccd1 _04451_
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10621_ _03395_ _03345_ _03411_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__o21ai_1
XFILLER_186_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__02435_ clknet_0__02435_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02435_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13340_ _05301_ vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__buf_4
XFILLER_194_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10552_ rbzero.debug_overlay.playerY\[2\] _03346_ rbzero.map_rom.a6 _03347_ vssd1
+ vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_168_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13271_ _06025_ _06027_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10483_ rbzero.tex_b0\[27\] rbzero.tex_b0\[26\] _03302_ vssd1 vssd1 vccd1 vccd1 _03308_
+ sky130_fd_sc_hd__mux2_1
XFILLER_154_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15010_ _07479_ _07697_ vssd1 vssd1 vccd1 vccd1 _07698_ sky130_fd_sc_hd__xnor2_2
X_12222_ _04970_ rbzero.wall_tracer.trackDistX\[-4\] _04971_ rbzero.wall_tracer.trackDistX\[-5\]
+ _04983_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__a221o_1
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12153_ _04913_ _04914_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__nand2_1
XFILLER_150_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11104_ rbzero.debug_overlay.playerY\[-3\] vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__inv_2
XFILLER_116_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16961_ _08862_ _08899_ _07961_ _08071_ vssd1 vssd1 vccd1 vccd1 _09567_ sky130_fd_sc_hd__or4_1
X_12084_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] vssd1
+ vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__nand2_1
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18700_ rbzero.debug_overlay.playerY\[-8\] _02588_ vssd1 vssd1 vccd1 vccd1 _02591_
+ sky130_fd_sc_hd__nor2_1
XFILLER_110_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19169__330 clknet_1_1__leaf__02748_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__inv_2
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15912_ rbzero.wall_tracer.trackDistX\[-8\] rbzero.wall_tracer.stepDistX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _08534_ sky130_fd_sc_hd__nand2_1
X_11035_ rbzero.row_render.size\[10\] rbzero.row_render.size\[9\] _03776_ _03820_
+ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__or4_4
X_19680_ clknet_leaf_80_i_clk _00611_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16892_ _09477_ _09498_ vssd1 vssd1 vccd1 vccd1 _09499_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18631_ _02534_ _02536_ _02537_ _02356_ vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__o211a_1
XFILLER_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15843_ _03395_ _08472_ vssd1 vssd1 vccd1 vccd1 _08473_ sky130_fd_sc_hd__nand2_1
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18562_ rbzero.pov.spi_buffer\[49\] rbzero.pov.spi_buffer\[50\] _02499_ vssd1 vssd1
+ vccd1 vccd1 _02500_ sky130_fd_sc_hd__mux2_1
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ _05505_ _05610_ _05741_ _05742_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__a2bb2o_1
X_15774_ _03469_ _08443_ _08446_ vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__o21a_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17513_ _01792_ _01790_ _01777_ vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__o21ai_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ _07412_ _07067_ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__nor2_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18493_ _02463_ vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__clkbuf_1
X_11937_ net69 _04665_ _04669_ _03910_ _04711_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__a221o_1
XFILLER_75_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _01735_ _01736_ _01738_ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__o21ai_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11868_ net13 _04638_ _04643_ _04632_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_21_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14656_ _07091_ _07156_ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__nor2_1
X_10819_ _03567_ _03603_ _03604_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__or3_1
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13607_ _06173_ _06316_ _06315_ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__nand3_1
X_17375_ rbzero.debug_overlay.playerX\[0\] _03373_ _09620_ vssd1 vssd1 vccd1 vccd1
+ _01680_ sky130_fd_sc_hd__mux2_1
X_14587_ _06940_ _07024_ _07037_ _06969_ vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__o22a_1
XFILLER_14_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11799_ net40 _04569_ _04570_ _03537_ _04575_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__a221o_1
XFILLER_13_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16326_ _08908_ _08937_ vssd1 vssd1 vccd1 vccd1 _08938_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13538_ _06293_ _06287_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__xor2_1
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16257_ _08107_ _08081_ vssd1 vssd1 vccd1 vccd1 _08869_ sky130_fd_sc_hd__nor2_1
X_13469_ _06208_ _06225_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__nor2_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15208_ _06853_ _07893_ _07894_ _07161_ vssd1 vssd1 vccd1 vccd1 _07895_ sky130_fd_sc_hd__o31a_1
X_16188_ _08392_ _08799_ _08800_ vssd1 vssd1 vccd1 vccd1 _08801_ sky130_fd_sc_hd__o21ai_1
XFILLER_142_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15139_ _07826_ _04929_ _06851_ vssd1 vssd1 vccd1 vccd1 _07827_ sky130_fd_sc_hd__mux2_2
XFILLER_114_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19947_ net176 _00878_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19878_ clknet_leaf_22_i_clk _00809_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18829_ rbzero.debug_overlay.vplaneX\[-2\] _02634_ vssd1 vssd1 vccd1 vccd1 _02677_
+ sky130_fd_sc_hd__and2_1
XFILLER_96_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18909__96 clknet_1_0__leaf__02441_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__inv_2
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20018_ clknet_leaf_92_i_clk _00949_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09829_ rbzero.tex_r1\[15\] rbzero.tex_r1\[16\] _02954_ vssd1 vssd1 vccd1 vccd1 _02963_
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12840_ _05589_ _05596_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _05527_ _05471_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__nor2_1
XFILLER_15_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ gpout0.vpos\[1\] vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__buf_2
X_14510_ _07154_ vssd1 vssd1 vccd1 vccd1 _07198_ sky130_fd_sc_hd__clkbuf_4
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ rbzero.debug_overlay.playerY\[-3\] rbzero.debug_overlay.playerX\[-3\] _06851_
+ vssd1 vssd1 vccd1 vccd1 _08175_ sky130_fd_sc_hd__mux2_1
XFILLER_159_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11653_ rbzero.tex_b1\[29\] rbzero.tex_b1\[28\] _04376_ vssd1 vssd1 vccd1 vccd1 _04434_
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14441_ _06733_ _06738_ _07103_ vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__nand3_1
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10604_ _03343_ _03358_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__xnor2_1
X_17160_ _01497_ _01503_ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__xnor2_1
X_14372_ _07054_ _07059_ vssd1 vssd1 vccd1 vccd1 _07060_ sky130_fd_sc_hd__nor2_1
XFILLER_80_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11584_ rbzero.tex_b0\[10\] _03700_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__and2_1
XFILLER_70_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16111_ _08611_ _08612_ _08723_ vssd1 vssd1 vccd1 vccd1 _08724_ sky130_fd_sc_hd__o21a_1
X_13323_ _05990_ _06061_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__or2_1
X_10535_ rbzero.tex_b0\[2\] rbzero.tex_b0\[1\] _02983_ vssd1 vssd1 vccd1 vccd1 _03335_
+ sky130_fd_sc_hd__mux2_1
XFILLER_127_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17091_ _09595_ _09694_ _09695_ vssd1 vssd1 vccd1 vccd1 _09696_ sky130_fd_sc_hd__o21ba_1
XFILLER_122_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16042_ _08645_ _08655_ vssd1 vssd1 vccd1 vccd1 _08656_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13254_ _05953_ _06007_ _06010_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__o21a_1
X_10466_ rbzero.tex_b0\[35\] rbzero.tex_b0\[34\] _03291_ vssd1 vssd1 vccd1 vccd1 _03299_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12205_ rbzero.wall_tracer.trackDistY\[0\] _04966_ vssd1 vssd1 vccd1 vccd1 _04967_
+ sky130_fd_sc_hd__nand2_1
X_13185_ _05888_ _05908_ _05941_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__a21oi_2
XFILLER_151_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10397_ rbzero.tex_b1\[3\] rbzero.tex_b1\[4\] _03254_ vssd1 vssd1 vccd1 vccd1 _03263_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19801_ clknet_leaf_16_i_clk _00732_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12136_ _04859_ _04860_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__xnor2_2
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17993_ rbzero.pov.spi_buffer\[49\] rbzero.pov.ready_buffer\[49\] _02197_ vssd1 vssd1
+ vccd1 vccd1 _02198_ sky130_fd_sc_hd__mux2_1
X_19732_ clknet_leaf_93_i_clk _00663_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_16944_ _09021_ _09036_ vssd1 vssd1 vccd1 vccd1 _09550_ sky130_fd_sc_hd__nor2_1
XFILLER_150_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12067_ net72 rbzero.wall_tracer.state\[7\] _04834_ vssd1 vssd1 vccd1 vccd1 _04835_
+ sky130_fd_sc_hd__and3_1
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11018_ rbzero.row_render.size\[4\] _03773_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19663_ clknet_leaf_4_i_clk _00594_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_16875_ _09480_ _09481_ vssd1 vssd1 vccd1 vccd1 _09482_ sky130_fd_sc_hd__or2_1
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18614_ _02526_ vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15826_ _08460_ vssd1 vssd1 vccd1 vccd1 _08463_ sky130_fd_sc_hd__buf_4
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19594_ clknet_leaf_44_i_clk _00525_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18545_ rbzero.pov.spi_buffer\[41\] rbzero.pov.spi_buffer\[42\] _02488_ vssd1 vssd1
+ vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
XFILLER_52_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15757_ _02899_ _08438_ vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__nor2_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _05700_ _05725_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14708_ _06993_ _07048_ vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__nor2_1
XFILLER_166_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18476_ _02454_ vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__clkbuf_1
X_15688_ _08232_ _08233_ _08230_ vssd1 vssd1 vccd1 vccd1 _08371_ sky130_fd_sc_hd__o21a_1
XFILLER_60_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17427_ _01722_ _01723_ _01724_ _08460_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__a31o_1
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14639_ _07292_ _07317_ vssd1 vssd1 vccd1 vccd1 _07327_ sky130_fd_sc_hd__nor2_1
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17358_ _01671_ vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16309_ _08909_ _08919_ vssd1 vssd1 vccd1 vccd1 _08921_ sky130_fd_sc_hd__or2_1
X_17289_ rbzero.wall_tracer.trackDistY\[4\] rbzero.wall_tracer.stepDistY\[4\] vssd1
+ vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__or2_1
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19244__18 clknet_1_0__leaf__02755_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__inv_2
XFILLER_84_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10320_ rbzero.tex_b1\[40\] rbzero.tex_b1\[41\] _03221_ vssd1 vssd1 vccd1 vccd1 _03223_
+ sky130_fd_sc_hd__mux2_1
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20498_ clknet_leaf_41_i_clk _01429_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10251_ _03186_ vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19051__224 clknet_1_1__leaf__02736_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__inv_2
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10182_ _03150_ vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18428__68 clknet_1_1__leaf__02438_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__inv_2
XFILLER_120_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14990_ _07676_ _07677_ vssd1 vssd1 vccd1 vccd1 _07678_ sky130_fd_sc_hd__nand2_1
XFILLER_94_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13941_ _06664_ _06690_ _06691_ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__a21oi_1
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16660_ _09048_ _09050_ vssd1 vssd1 vccd1 vccd1 _09269_ sky130_fd_sc_hd__nand2_2
XFILLER_75_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13872_ _05272_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__clkbuf_4
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15611_ _08185_ _08293_ vssd1 vssd1 vccd1 vccd1 _08295_ sky130_fd_sc_hd__or2_1
XFILLER_90_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12823_ _05577_ _05579_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__or2_1
XFILLER_61_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16591_ _09082_ _09086_ vssd1 vssd1 vccd1 vccd1 _09201_ sky130_fd_sc_hd__nand2_1
XFILLER_188_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18330_ rbzero.spi_registers.spi_cmd\[3\] rbzero.spi_registers.spi_cmd\[2\] rbzero.spi_registers.spi_done
+ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__and3b_1
XFILLER_188_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15542_ _08097_ _08224_ _08225_ vssd1 vssd1 vccd1 vccd1 _08226_ sky130_fd_sc_hd__a21o_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12754_ _05500_ _05487_ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__xnor2_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _04477_ _04478_ _04484_ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__a21oi_1
X_18261_ rbzero.spi_registers.spi_buffer\[0\] rbzero.spi_registers.new_sky\[0\] _02361_
+ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__mux2_1
X_15473_ _08026_ _08027_ _08030_ _08031_ _08006_ vssd1 vssd1 vccd1 vccd1 _08158_ sky130_fd_sc_hd__a32oi_2
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _05414_ _05441_ _05209_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__o21a_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _01547_ _01548_ _01549_ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__o21ai_1
X_11636_ rbzero.tex_b1\[63\] rbzero.tex_b1\[62\] _03616_ vssd1 vssd1 vccd1 vccd1 _04417_
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14424_ _06849_ _04888_ vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__or2_1
X_18192_ rbzero.spi_registers.new_leak\[2\] _02310_ _02315_ _02314_ vssd1 vssd1 vccd1
+ vccd1 _00779_ sky130_fd_sc_hd__o211a_1
XFILLER_168_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17143_ _01483_ _01486_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__xnor2_1
XFILLER_155_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11567_ _03688_ _04323_ _04331_ _04348_ _03718_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__a311o_1
X_14355_ _03491_ rbzero.wall_tracer.stepDistY\[-9\] _06906_ vssd1 vssd1 vccd1 vccd1
+ _07043_ sky130_fd_sc_hd__a21oi_1
XFILLER_200_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10518_ _03326_ vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13306_ _06060_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__xnor2_1
X_17074_ _09677_ _09678_ vssd1 vssd1 vccd1 vccd1 _09679_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_1_1__f__02732_ clknet_0__02732_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02732_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_128_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14286_ _04890_ _05124_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__mux2_1
X_11498_ rbzero.tex_g1\[62\] _03925_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__and2_1
XFILLER_144_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16025_ _06875_ _07123_ vssd1 vssd1 vccd1 vccd1 _08639_ sky130_fd_sc_hd__or2_1
X_13237_ _05900_ _05905_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__xnor2_1
X_10449_ rbzero.tex_b0\[43\] rbzero.tex_b0\[42\] _03280_ vssd1 vssd1 vccd1 vccd1 _03290_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13168_ _05865_ _05866_ _05924_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__a21bo_1
XFILLER_152_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12119_ _04877_ _04878_ _04879_ _04880_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__o31a_1
X_13099_ _05687_ _05766_ _05852_ _05855_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__a2bb2o_1
X_17976_ rbzero.pov.spi_buffer\[41\] rbzero.pov.ready_buffer\[41\] _02186_ vssd1 vssd1
+ vccd1 vccd1 _02189_ sky130_fd_sc_hd__mux2_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19715_ clknet_leaf_3_i_clk _00646_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16927_ _09377_ _09381_ vssd1 vssd1 vccd1 vccd1 _09533_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_62_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19646_ clknet_leaf_46_i_clk _00577_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16858_ _09377_ _09382_ vssd1 vssd1 vccd1 vccd1 _09465_ sky130_fd_sc_hd__nand2_1
XFILLER_168_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15809_ rbzero.traced_texa\[-8\] _08457_ _08459_ rbzero.wall_tracer.visualWallDist\[-8\]
+ vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__a22o_1
X_19577_ clknet_leaf_33_i_clk _00508_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16789_ _09289_ _09291_ vssd1 vssd1 vccd1 vccd1 _09397_ sky130_fd_sc_hd__nor2_1
XFILLER_92_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_77_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18528_ rbzero.pov.spi_buffer\[33\] rbzero.pov.spi_buffer\[34\] _02477_ vssd1 vssd1
+ vccd1 vccd1 _02482_ sky130_fd_sc_hd__mux2_1
XFILLER_179_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18459_ rbzero.pov.spi_buffer\[0\] rbzero.pov.spi_buffer\[1\] _02444_ vssd1 vssd1
+ vccd1 vccd1 _02446_ sky130_fd_sc_hd__mux2_1
XFILLER_21_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20421_ net481 _01352_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20352_ net412 _01283_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19000__178 clknet_1_1__leaf__02731_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__inv_2
XFILLER_135_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20283_ net343 _01214_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__02752_ clknet_0__02752_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02752_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12470_ _05199_ _05132_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__nand2_2
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11421_ _03917_ _04202_ _04204_ _03689_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__o211a_1
XFILLER_138_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14140_ rbzero.wall_tracer.stepDistX\[7\] _06772_ _06825_ vssd1 vssd1 vccd1 vccd1
+ _06835_ sky130_fd_sc_hd__mux2_1
XFILLER_165_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11352_ rbzero.debug_overlay.playerY\[-2\] _04056_ _04084_ rbzero.debug_overlay.playerY\[-6\]
+ _04136_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__a221o_1
XFILLER_193_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10303_ rbzero.tex_b1\[48\] rbzero.tex_b1\[49\] _03210_ vssd1 vssd1 vccd1 vccd1 _03214_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14071_ rbzero.wall_tracer.visualWallDist\[-4\] _06796_ _06791_ rbzero.wall_tracer.trackDistX\[-4\]
+ _06797_ vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__o221a_1
X_11283_ _04051_ _04067_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__nor2_1
XFILLER_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13022_ _05473_ _05536_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__nor2_1
X_10234_ rbzero.tex_g0\[18\] rbzero.tex_g0\[17\] _03177_ vssd1 vssd1 vccd1 vccd1 _03178_
+ sky130_fd_sc_hd__mux2_1
X_18916__102 clknet_1_0__leaf__02723_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__inv_2
XFILLER_4_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17830_ _02090_ _02092_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__xnor2_1
X_10165_ rbzero.tex_g0\[50\] rbzero.tex_g0\[49\] _03132_ vssd1 vssd1 vccd1 vccd1 _03141_
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17761_ rbzero.debug_overlay.vplaneX\[-1\] _04100_ vssd1 vssd1 vccd1 vccd1 _02029_
+ sky130_fd_sc_hd__nor2_1
X_10096_ rbzero.tex_g1\[18\] rbzero.tex_g1\[19\] _03095_ vssd1 vssd1 vccd1 vccd1 _03105_
+ sky130_fd_sc_hd__mux2_1
X_14973_ _07617_ vssd1 vssd1 vccd1 vccd1 _07661_ sky130_fd_sc_hd__buf_2
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19500_ clknet_leaf_46_i_clk _00446_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[7\]
+ sky130_fd_sc_hd__dfxtp_4
X_16712_ _09318_ _09319_ vssd1 vssd1 vccd1 vccd1 _09320_ sky130_fd_sc_hd__nor2_1
X_13924_ _06610_ _06676_ _06664_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__mux2_1
X_17692_ _01961_ _01962_ _01964_ vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__nand3_1
XFILLER_75_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19431_ _01919_ _01928_ _01927_ _08464_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__a31o_1
XFILLER_74_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16643_ _09250_ _09251_ vssd1 vssd1 vccd1 vccd1 _09252_ sky130_fd_sc_hd__xnor2_1
X_13855_ _05349_ _06611_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__nor2_1
XFILLER_90_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12806_ _05392_ _05535_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__or2_1
X_19362_ _02839_ _02842_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__xnor2_1
X_16574_ _09181_ _09182_ vssd1 vssd1 vccd1 vccd1 _09184_ sky130_fd_sc_hd__nand2_1
XFILLER_34_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13786_ _06530_ _06541_ _06542_ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__o21bai_1
X_10998_ rbzero.row_render.size\[1\] _03499_ _03500_ rbzero.row_render.size\[0\] vssd1
+ vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__a211o_1
XFILLER_90_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18313_ rbzero.spi_registers.new_other\[2\] rbzero.spi_registers.spi_buffer\[2\]
+ _02388_ vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__mux2_1
X_18962__144 clknet_1_1__leaf__02727_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__inv_2
X_15525_ _07856_ _08081_ vssd1 vssd1 vccd1 vccd1 _08209_ sky130_fd_sc_hd__nor2_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12737_ _05210_ _05445_ _05446_ _05323_ _05448_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__a32o_4
X_19293_ rbzero.texV\[-6\] _02675_ _02709_ _02784_ vssd1 vssd1 vccd1 vccd1 _01411_
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ rbzero.spi_registers.vshift\[1\] _02349_ vssd1 vssd1 vccd1 vccd1 _02351_
+ sky130_fd_sc_hd__or2_1
XFILLER_30_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15456_ _08139_ _08140_ _07161_ vssd1 vssd1 vccd1 vccd1 _08141_ sky130_fd_sc_hd__o21ai_2
X_12668_ _05416_ _05417_ _05424_ _05209_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__nand4b_4
XFILLER_175_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14407_ _07078_ _06968_ _07094_ vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__or3_1
X_11619_ rbzero.tex_b1\[43\] rbzero.tex_b1\[42\] _03662_ vssd1 vssd1 vccd1 vccd1 _04400_
+ sky130_fd_sc_hd__mux2_1
XFILLER_129_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18175_ rbzero.spi_registers.new_mapd\[9\] _02289_ _02305_ _02301_ vssd1 vssd1 vccd1
+ vccd1 _00772_ sky130_fd_sc_hd__o211a_1
X_15387_ _07011_ _07269_ _07961_ _08071_ vssd1 vssd1 vccd1 vccd1 _08072_ sky130_fd_sc_hd__nor4_1
XFILLER_184_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12599_ _05274_ _05320_ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__xnor2_4
XFILLER_129_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17126_ _09133_ _09110_ _09676_ _01469_ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__o31a_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14338_ rbzero.debug_overlay.playerY\[-1\] rbzero.debug_overlay.playerY\[-2\] _06980_
+ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__or3_4
XFILLER_116_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17057_ _08896_ _08071_ vssd1 vssd1 vccd1 vccd1 _09662_ sky130_fd_sc_hd__or2_1
X_14269_ rbzero.debug_overlay.playerY\[-5\] _06922_ rbzero.debug_overlay.playerY\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__o21ai_1
XFILLER_143_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16008_ _07865_ _08081_ vssd1 vssd1 vccd1 vccd1 _08622_ sky130_fd_sc_hd__nor2_1
XFILLER_143_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__02746_ _02746_ vssd1 vssd1 vccd1 vccd1 clknet_0__02746_ sky130_fd_sc_hd__clkbuf_16
XFILLER_171_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ rbzero.pov.spi_buffer\[33\] rbzero.pov.ready_buffer\[33\] _02175_ vssd1 vssd1
+ vccd1 vccd1 _02180_ sky130_fd_sc_hd__mux2_1
XFILLER_100_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18407__49 clknet_1_0__leaf__02436_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__inv_2
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19629_ clknet_leaf_53_i_clk _00560_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19080__250 clknet_1_0__leaf__02739_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__inv_2
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20404_ net464 _01335_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20335_ net395 _01266_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_122_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20266_ net326 _01197_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 o_gpout[5] sky130_fd_sc_hd__clkbuf_1
XFILLER_143_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20197_ net257 _01128_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_49_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ net53 _04730_ _04724_ net50 vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__a22o_1
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10921_ rbzero.tex_r0\[27\] rbzero.tex_r0\[26\] _03649_ vssd1 vssd1 vccd1 vccd1 _03707_
+ sky130_fd_sc_hd__mux2_1
X_19163__325 clknet_1_1__leaf__02747_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__inv_2
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__02735_ clknet_0__02735_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02735_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10852_ _03636_ _03637_ rbzero.row_render.wall\[1\] vssd1 vssd1 vccd1 vccd1 _03638_
+ sky130_fd_sc_hd__a21bo_1
X_13640_ _06231_ _06396_ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__nor2_1
XFILLER_71_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ rbzero.traced_texVinit\[10\] rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 _03569_
+ sky130_fd_sc_hd__xor2_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _06305_ _06326_ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__nor2_1
XFILLER_52_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ _07530_ _07138_ _07137_ _07581_ vssd1 vssd1 vccd1 vccd1 _07996_ sky130_fd_sc_hd__o22a_1
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _05238_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__inv_2
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16290_ _08898_ _08900_ vssd1 vssd1 vccd1 vccd1 _08902_ sky130_fd_sc_hd__and2_1
XFILLER_13_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15241_ _07832_ _07927_ vssd1 vssd1 vccd1 vccd1 _07928_ sky130_fd_sc_hd__xnor2_2
XFILLER_200_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12453_ _05209_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__buf_4
XFILLER_184_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11404_ _03614_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__clkbuf_8
XFILLER_166_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15172_ _07855_ _07858_ vssd1 vssd1 vccd1 vccd1 _07859_ sky130_fd_sc_hd__xnor2_1
X_12384_ _05056_ _05030_ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__or2b_2
XFILLER_181_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11335_ rbzero.debug_overlay.facingX\[-4\] _04089_ _04090_ rbzero.debug_overlay.facingX\[-8\]
+ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__a22o_1
X_14123_ _06826_ vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__clkbuf_1
X_19980_ net209 _00911_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11266_ _04035_ _04050_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__nand2_4
X_14054_ _06787_ _03496_ _06788_ rbzero.wall_tracer.trackDistX\[-11\] _03485_ vssd1
+ vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__o221a_1
XFILLER_140_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10217_ rbzero.tex_g0\[26\] rbzero.tex_g0\[25\] _03166_ vssd1 vssd1 vccd1 vccd1 _03169_
+ sky130_fd_sc_hd__mux2_1
X_13005_ _05700_ _05725_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__and2_1
X_18862_ _03852_ _04503_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__nor2_1
X_11197_ rbzero.tex_r1\[27\] _03936_ _03981_ _03726_ vssd1 vssd1 vccd1 vccd1 _03982_
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17813_ _02000_ rbzero.wall_tracer.rayAddendX\[8\] vssd1 vssd1 vccd1 vccd1 _02077_
+ sky130_fd_sc_hd__xnor2_1
X_10148_ _02983_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__clkbuf_4
X_18793_ rbzero.pov.ready_buffer\[24\] _02644_ _02656_ _02651_ vssd1 vssd1 vccd1 vccd1
+ _01039_ sky130_fd_sc_hd__a211o_1
X_17744_ _01985_ rbzero.wall_tracer.rayAddendX\[3\] vssd1 vssd1 vccd1 vccd1 _02013_
+ sky130_fd_sc_hd__nor2_1
X_10079_ _03096_ vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__clkbuf_1
X_14956_ _07630_ _07633_ vssd1 vssd1 vccd1 vccd1 _07644_ sky130_fd_sc_hd__or2_1
XFILLER_48_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13907_ _06603_ _06633_ _06660_ _05271_ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__a211o_1
X_17675_ _01722_ _01948_ _01949_ _08460_ vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__a31o_1
X_14887_ _07544_ _07568_ vssd1 vssd1 vccd1 vccd1 _07575_ sky130_fd_sc_hd__xor2_1
XFILLER_36_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19414_ _01705_ _02874_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16626_ _08888_ _09110_ vssd1 vssd1 vccd1 vccd1 _09235_ sky130_fd_sc_hd__nor2_1
XFILLER_63_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13838_ _06575_ _06586_ _06593_ _06594_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__a31o_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19345_ rbzero.traced_texa\[3\] rbzero.texV\[3\] vssd1 vssd1 vccd1 vccd1 _02828_
+ sky130_fd_sc_hd__or2_1
X_16557_ _09050_ _09166_ vssd1 vssd1 vccd1 vccd1 _09167_ sky130_fd_sc_hd__and2_1
XFILLER_50_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13769_ _06514_ _06525_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__and2b_1
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15508_ _07011_ _08191_ vssd1 vssd1 vccd1 vccd1 _08192_ sky130_fd_sc_hd__or2_1
X_19276_ _02767_ _02770_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__xnor2_1
X_16488_ _08985_ _09000_ _08998_ vssd1 vssd1 vccd1 vccd1 _09098_ sky130_fd_sc_hd__a21o_1
XFILLER_175_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18227_ _02339_ vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15439_ _08122_ _08123_ vssd1 vssd1 vccd1 vccd1 _08124_ sky130_fd_sc_hd__nand2_1
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18158_ rbzero.spi_registers.new_mapd\[13\] _02290_ _02296_ _02275_ vssd1 vssd1 vccd1
+ vccd1 _00764_ sky130_fd_sc_hd__o211a_1
XFILLER_141_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17109_ _09710_ _09711_ _09712_ _04946_ vssd1 vssd1 vccd1 vccd1 _09714_ sky130_fd_sc_hd__a31o_1
XFILLER_117_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18089_ _02249_ vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20120_ clknet_leaf_91_i_clk _01051_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-6\]
+ sky130_fd_sc_hd__dfxtp_2
X_09931_ _03018_ vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__02729_ _02729_ vssd1 vssd1 vccd1 vccd1 clknet_0__02729_ sky130_fd_sc_hd__clkbuf_16
X_20051_ clknet_leaf_82_i_clk _00982_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[67\]
+ sky130_fd_sc_hd__dfxtp_1
X_09862_ _02980_ vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__clkbuf_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19112__279 clknet_1_0__leaf__02742_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__inv_2
X_09793_ _02944_ vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19006__184 clknet_1_0__leaf__02731_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__inv_2
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11120_ gpout0.vpos\[8\] vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__clkbuf_4
XFILLER_107_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20318_ net378 _01249_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18991__170 clknet_1_1__leaf__02730_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__inv_2
X_11051_ _03832_ _03833_ _03836_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__or3b_1
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20249_ net309 _01180_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10002_ _03055_ vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14810_ _07463_ _07465_ vssd1 vssd1 vccd1 vccd1 _07498_ sky130_fd_sc_hd__xnor2_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ rbzero.row_render.size\[4\] _08456_ _06705_ _08455_ vssd1 vssd1 vccd1 vccd1
+ _00496_ sky130_fd_sc_hd__a22o_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14741_ _06932_ _06978_ vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__or2_1
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ _03459_ _03469_ net27 vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__mux2_1
Xtop_ew_algofoogle_105 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_105/HI zeros[14]
+ sky130_fd_sc_hd__conb_1
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_116 vssd1 vssd1 vccd1 vccd1 ones[9] top_ew_algofoogle_116/LO sky130_fd_sc_hd__conb_1
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10904_ _03615_ vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__clkbuf_8
X_17460_ rbzero.wall_tracer.rayAddendY\[-1\] _08447_ _01754_ _01714_ vssd1 vssd1 vccd1
+ vccd1 _01755_ sky130_fd_sc_hd__a22o_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _07073_ _07064_ vssd1 vssd1 vccd1 vccd1 _07360_ sky130_fd_sc_hd__xnor2_1
X_11884_ net43 _04626_ _04627_ _03911_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__a22o_1
XFILLER_33_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16411_ _09021_ _08896_ _08893_ _08892_ vssd1 vssd1 vccd1 vccd1 _09022_ sky130_fd_sc_hd__o31a_1
X_13623_ _06357_ _06378_ _06379_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__a21oi_1
X_10835_ rbzero.row_render.texu\[0\] _03620_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__nor2_1
XFILLER_73_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17391_ _01692_ vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16342_ _08952_ _08953_ vssd1 vssd1 vccd1 vccd1 _08954_ sky130_fd_sc_hd__xnor2_4
XFILLER_198_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13554_ _06103_ _05992_ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__nor2_1
XFILLER_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10766_ rbzero.texV\[3\] _03551_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__xor2_1
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12505_ _05238_ _05242_ _05261_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__or3_1
X_16273_ _06858_ _08252_ vssd1 vssd1 vccd1 vccd1 _08885_ sky130_fd_sc_hd__nor2_1
XFILLER_146_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13485_ _06008_ _05995_ _06151_ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__o21bai_1
X_10697_ rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__buf_2
XFILLER_186_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18012_ _02207_ vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__clkbuf_1
X_15224_ _07764_ _07769_ vssd1 vssd1 vccd1 vccd1 _07911_ sky130_fd_sc_hd__nor2_1
XFILLER_126_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12436_ _05189_ _05192_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__or2b_1
XFILLER_201_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15155_ _07709_ _07834_ _07841_ vssd1 vssd1 vccd1 vccd1 _07842_ sky130_fd_sc_hd__and3_1
XFILLER_126_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12367_ _05121_ _05123_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__xnor2_2
XFILLER_181_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14106_ _06817_ vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__clkbuf_1
X_11318_ rbzero.debug_overlay.vplaneX\[-9\] _04081_ _04089_ _04102_ vssd1 vssd1 vccd1
+ vccd1 _04103_ sky130_fd_sc_hd__a22o_1
X_19963_ net192 _00894_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[43\] sky130_fd_sc_hd__dfxtp_1
X_15086_ _07771_ _07772_ vssd1 vssd1 vccd1 vccd1 _07774_ sky130_fd_sc_hd__nand2_1
X_12298_ rbzero.debug_overlay.facingX\[0\] rbzero.wall_tracer.rayAddendX\[8\] vssd1
+ vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__and2_1
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14037_ _05395_ _06634_ _05373_ vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__a21oi_1
X_11249_ _03476_ _04033_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__and2_2
XFILLER_80_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19894_ clknet_leaf_18_i_clk _00825_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_95_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18845_ rbzero.debug_overlay.vplaneY\[-5\] _02634_ vssd1 vssd1 vccd1 vccd1 _02685_
+ sky130_fd_sc_hd__and2_1
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18776_ rbzero.pov.ready_buffer\[38\] _02644_ _02647_ _02559_ vssd1 vssd1 vccd1 vccd1
+ _01031_ sky130_fd_sc_hd__a211o_1
X_15988_ _08352_ _08599_ _08600_ vssd1 vssd1 vccd1 vccd1 _08602_ sky130_fd_sc_hd__and3_1
XFILLER_67_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17727_ _01980_ _01995_ _01991_ vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__or3_1
XFILLER_76_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14939_ _07622_ _07626_ vssd1 vssd1 vccd1 vccd1 _07627_ sky130_fd_sc_hd__nand2_1
XFILLER_82_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18397__40 clknet_1_0__leaf__02435_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__inv_2
XFILLER_35_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17658_ _04102_ rbzero.wall_tracer.rayAddendX\[-4\] vssd1 vssd1 vccd1 vccd1 _01934_
+ sky130_fd_sc_hd__nand2_1
XFILLER_169_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16609_ _07993_ _07960_ _08071_ _08643_ vssd1 vssd1 vccd1 vccd1 _09218_ sky130_fd_sc_hd__o22a_1
XFILLER_51_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17589_ _01862_ _01870_ _01874_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__a21o_1
XFILLER_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19328_ _02813_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__inv_2
XFILLER_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19259_ gpout5.clk_div\[1\] gpout5.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__or2_1
XFILLER_192_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19192__351 clknet_1_1__leaf__02750_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__inv_2
XFILLER_176_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20103_ clknet_leaf_88_i_clk _01034_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
X_09914_ _03009_ vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20034_ clknet_leaf_7_i_clk _00965_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_09845_ _02971_ vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__clkbuf_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ _02935_ vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__clkbuf_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10620_ _03395_ _03345_ _03375_ _03354_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__a22o_1
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__02434_ clknet_0__02434_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02434_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_195_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10551_ rbzero.debug_overlay.playerY\[3\] vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__inv_2
XFILLER_195_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10482_ _03307_ vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__clkbuf_1
X_13270_ _05961_ _05968_ _06026_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__a21oi_1
XFILLER_194_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12221_ _04971_ rbzero.wall_tracer.trackDistX\[-5\] _04972_ rbzero.wall_tracer.trackDistX\[-6\]
+ _04982_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__o221a_1
XFILLER_151_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12152_ _04870_ _04873_ _04912_ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__or3b_1
XFILLER_68_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11103_ gpout0.vpos\[1\] rbzero.debug_overlay.playerY\[-2\] vssd1 vssd1 vccd1 vccd1
+ _03889_ sky130_fd_sc_hd__xnor2_1
X_16960_ _08899_ _07961_ vssd1 vssd1 vccd1 vccd1 _09566_ sky130_fd_sc_hd__nor2_1
X_12083_ _04843_ _04844_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__nand2_1
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15911_ rbzero.wall_tracer.trackDistX\[-8\] rbzero.wall_tracer.stepDistX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _08533_ sky130_fd_sc_hd__or2_1
X_11034_ _03792_ _03795_ _03818_ _03819_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_104_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16891_ _09496_ _09497_ vssd1 vssd1 vccd1 vccd1 _09498_ sky130_fd_sc_hd__nand2_1
XFILLER_76_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18630_ _07145_ _02533_ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__nand2_1
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15842_ _03362_ _06914_ vssd1 vssd1 vccd1 vccd1 _08472_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18561_ _02443_ vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__clkbuf_4
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _03469_ _08443_ _08438_ vssd1 vssd1 vccd1 vccd1 _08446_ sky130_fd_sc_hd__a21oi_1
X_12985_ _05484_ _05473_ _05505_ _05425_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__o211a_1
XFILLER_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ _01790_ _01793_ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__nand2_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _07068_ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__inv_2
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18492_ rbzero.pov.spi_buffer\[16\] rbzero.pov.spi_buffer\[17\] _02455_ vssd1 vssd1
+ vccd1 vccd1 _02463_ sky130_fd_sc_hd__mux2_1
X_11936_ net47 _04668_ _04710_ _04666_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__a22o_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17443_ _01735_ _01736_ _01738_ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__or3_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14655_ _07297_ _07298_ vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__xnor2_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _04639_ _04623_ _04640_ _04635_ _04642_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__a32o_2
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13606_ _06362_ _06340_ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__xnor2_1
X_10818_ _03566_ _03550_ _03558_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__nor3_1
XFILLER_14_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17374_ _01679_ vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14586_ _06940_ _07273_ _07247_ vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__or3_1
X_11798_ net49 _04566_ _04568_ net39 vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a22o_1
XFILLER_13_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16325_ _08935_ _08936_ vssd1 vssd1 vccd1 vccd1 _08937_ sky130_fd_sc_hd__nor2_1
X_13537_ _06287_ _06293_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__or2b_1
XFILLER_9_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10749_ _02902_ _03467_ gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__a21oi_4
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16256_ _08866_ _08867_ vssd1 vssd1 vccd1 vccd1 _08868_ sky130_fd_sc_hd__nand2_1
XFILLER_173_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13468_ _06222_ _06223_ vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__and2_1
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15207_ _06759_ _06764_ _07165_ _06767_ vssd1 vssd1 vccd1 vccd1 _07894_ sky130_fd_sc_hd__o31a_1
X_12419_ _05155_ _05156_ _05161_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__o21a_1
X_16187_ _07661_ _08391_ _08678_ _07662_ vssd1 vssd1 vccd1 vccd1 _08800_ sky130_fd_sc_hd__o22ai_1
XFILLER_126_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13399_ _06155_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__clkbuf_4
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15138_ _07825_ vssd1 vssd1 vccd1 vccd1 _07826_ sky130_fd_sc_hd__clkbuf_4
XFILLER_142_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19946_ net175 _00877_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[26\] sky130_fd_sc_hd__dfxtp_1
X_15069_ _07754_ vssd1 vssd1 vccd1 vccd1 _07757_ sky130_fd_sc_hd__buf_2
XFILLER_114_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19877_ clknet_leaf_21_i_clk _00808_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_sky
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18828_ rbzero.pov.ready_buffer\[17\] _02663_ _02676_ _02672_ vssd1 vssd1 vccd1 vccd1
+ _01054_ sky130_fd_sc_hd__o211a_1
XFILLER_67_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18759_ _02635_ vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__buf_2
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19118__285 clknet_1_1__leaf__02742_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__inv_2
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20017_ clknet_leaf_92_i_clk _00948_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09828_ _02962_ vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09759_ _02926_ vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _05526_ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__clkbuf_4
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ gpout0.vpos\[0\] vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__buf_2
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _07086_ _07127_ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__xnor2_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _03688_ _04415_ _04432_ _03719_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__o211a_1
X_19199__357 clknet_1_0__leaf__02751_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__inv_2
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10603_ rbzero.map_rom.f2 rbzero.map_rom.b6 vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__or2_1
X_18391__35 clknet_1_1__leaf__02434_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__inv_2
X_14371_ _07055_ _07058_ _07056_ vssd1 vssd1 vccd1 vccd1 _07059_ sky130_fd_sc_hd__a21oi_1
X_11583_ _03671_ _04360_ _04364_ _03679_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__a211o_1
XFILLER_22_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16110_ _08613_ _08614_ vssd1 vssd1 vccd1 vccd1 _08723_ sky130_fd_sc_hd__or2b_1
XFILLER_155_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13322_ _06000_ _06067_ _06078_ vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__o21ai_1
XFILLER_196_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17090_ _09575_ _09576_ _09573_ vssd1 vssd1 vccd1 vccd1 _09695_ sky130_fd_sc_hd__a21oi_1
X_10534_ _03334_ vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16041_ _08653_ _08654_ vssd1 vssd1 vccd1 vccd1 _08655_ sky130_fd_sc_hd__nor2_1
X_10465_ _03298_ vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__clkbuf_1
X_13253_ _05235_ _05616_ _05954_ _06009_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__a31oi_1
XFILLER_171_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12204_ rbzero.wall_tracer.trackDistX\[0\] vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__inv_2
XFILLER_108_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10396_ _03262_ vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13184_ _05939_ _05940_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__nand2_1
XFILLER_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19800_ clknet_leaf_16_i_clk _00731_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12135_ rbzero.wall_tracer.rayAddendY\[-3\] rbzero.wall_tracer.rayAddendY\[-2\] _04894_
+ _04896_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__or4bb_1
XFILLER_2_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17992_ _02141_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__clkbuf_4
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16943_ _09485_ _09546_ _09548_ vssd1 vssd1 vccd1 vccd1 _09549_ sky130_fd_sc_hd__a21oi_1
X_19731_ clknet_leaf_94_i_clk _00662_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12066_ _04827_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__buf_6
XFILLER_96_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11017_ _03774_ _03802_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__nand2_1
X_16874_ _09007_ _09256_ _09039_ _09009_ vssd1 vssd1 vccd1 vccd1 _09481_ sky130_fd_sc_hd__o22a_1
X_19662_ clknet_leaf_4_i_clk _00593_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18613_ rbzero.pov.mosi rbzero.pov.mosi_buffer\[0\] _04827_ vssd1 vssd1 vccd1 vccd1
+ _02526_ sky130_fd_sc_hd__mux2_1
XFILLER_49_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15825_ rbzero.traced_texa\[5\] _08461_ _08462_ rbzero.wall_tracer.visualWallDist\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__a22o_1
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19593_ clknet_leaf_40_i_clk _00524_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18544_ _02490_ vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__clkbuf_1
X_15756_ _08437_ vssd1 vssd1 vccd1 vccd1 _08438_ sky130_fd_sc_hd__clkbuf_2
XFILLER_18_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12968_ _05722_ _05724_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__xor2_1
XFILLER_92_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14707_ _06998_ _07394_ vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__or2_1
XFILLER_166_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18475_ rbzero.pov.spi_buffer\[8\] rbzero.pov.spi_buffer\[9\] _02444_ vssd1 vssd1
+ vccd1 vccd1 _02454_ sky130_fd_sc_hd__mux2_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11919_ _04503_ _04672_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__nor2_1
X_15687_ _08365_ _08369_ vssd1 vssd1 vccd1 vccd1 _08370_ sky130_fd_sc_hd__xor2_1
XFILLER_61_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ _05467_ _05483_ _05505_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__a21o_1
XFILLER_61_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__nand2_1
X_14638_ _07319_ _07325_ vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17357_ rbzero.spi_registers.new_mapd\[7\] rbzero.spi_registers.spi_buffer\[7\] _01663_
+ vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__mux2_1
XFILLER_158_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14569_ rbzero.wall_tracer.visualWallDist\[3\] _07256_ vssd1 vssd1 vccd1 vccd1 _07257_
+ sky130_fd_sc_hd__nand2_1
XFILLER_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16308_ _08909_ _08919_ vssd1 vssd1 vccd1 vccd1 _08920_ sky130_fd_sc_hd__nand2_1
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17288_ rbzero.wall_tracer.trackDistY\[4\] rbzero.wall_tracer.stepDistY\[4\] vssd1
+ vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__nand2_1
X_16239_ _08850_ vssd1 vssd1 vccd1 vccd1 _08851_ sky130_fd_sc_hd__inv_2
XFILLER_146_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19929_ net158 _00860_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20497_ clknet_leaf_37_i_clk _01428_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_164_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10250_ rbzero.tex_g0\[10\] rbzero.tex_g0\[9\] _03177_ vssd1 vssd1 vccd1 vccd1 _03186_
+ sky130_fd_sc_hd__mux2_1
XFILLER_106_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10181_ rbzero.tex_g0\[43\] rbzero.tex_g0\[42\] _03144_ vssd1 vssd1 vccd1 vccd1 _03150_
+ sky130_fd_sc_hd__mux2_1
XFILLER_191_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13940_ _06664_ _06676_ vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__nor2_1
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13871_ _05410_ _06613_ _06627_ _05333_ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__a211o_1
XFILLER_189_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15610_ _08185_ _08293_ vssd1 vssd1 vccd1 vccd1 _08294_ sky130_fd_sc_hd__nand2_2
XFILLER_62_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12822_ _05548_ _05578_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16590_ _09198_ _09199_ vssd1 vssd1 vccd1 vccd1 _09200_ sky130_fd_sc_hd__nand2_1
XFILLER_90_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15541_ _06858_ _07735_ _07097_ _06875_ vssd1 vssd1 vccd1 vccd1 _08225_ sky130_fd_sc_hd__o22a_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12753_ _05485_ _05504_ _05506_ _05509_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__a22oi_2
XFILLER_43_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ _02360_ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__clkbuf_4
X_11704_ _03499_ _04479_ _04482_ _04020_ _04483_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__o2111a_1
X_15472_ _08128_ _08156_ vssd1 vssd1 vccd1 vccd1 _08157_ sky130_fd_sc_hd__xnor2_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12684_ _05440_ _05345_ _05329_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__mux2_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _01547_ _01548_ _01549_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__or3_1
X_14423_ _06717_ _06726_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__xnor2_1
X_11635_ rbzero.tex_b1\[61\] rbzero.tex_b1\[60\] _03616_ vssd1 vssd1 vccd1 vccd1 _04416_
+ sky130_fd_sc_hd__mux2_1
X_18191_ rbzero.floor_leak\[2\] _02311_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__or2_1
XFILLER_129_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17142_ _09637_ _01485_ vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14354_ _07025_ _07038_ _07041_ vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__a21bo_1
XFILLER_129_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11566_ _03704_ _04335_ _04339_ _04347_ _03684_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__o311a_1
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13305_ _06001_ _06061_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__nor2_1
XFILLER_116_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__02731_ clknet_0__02731_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02731_
+ sky130_fd_sc_hd__clkbuf_16
X_17073_ _09133_ _09110_ vssd1 vssd1 vccd1 vccd1 _09678_ sky130_fd_sc_hd__nor2_1
X_10517_ rbzero.tex_b0\[11\] rbzero.tex_b0\[10\] _03324_ vssd1 vssd1 vccd1 vccd1 _03326_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14285_ _03490_ rbzero.wall_tracer.stepDistY\[-7\] _04947_ vssd1 vssd1 vccd1 vccd1
+ _06973_ sky130_fd_sc_hd__a21oi_1
X_11497_ _04276_ _04279_ _03671_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__mux2_1
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16024_ _08379_ _08384_ vssd1 vssd1 vccd1 vccd1 _08638_ sky130_fd_sc_hd__nand2_1
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13236_ _05990_ _05992_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__nor2_1
XFILLER_196_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10448_ _03289_ vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13167_ _05867_ _05868_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__or2b_1
XFILLER_3_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10379_ _03253_ vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12118_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[10\] vssd1
+ vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__nand2_1
XFILLER_111_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17975_ _02188_ vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__clkbuf_1
X_13098_ _05687_ _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19714_ clknet_leaf_2_i_clk _00645_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16926_ _09283_ _09471_ _09280_ vssd1 vssd1 vccd1 vccd1 _09532_ sky130_fd_sc_hd__a21bo_1
X_12049_ clknet_leaf_27_i_clk _04794_ _04791_ _04821_ net35 vssd1 vssd1 vccd1 vccd1
+ _04822_ sky130_fd_sc_hd__a2111oi_2
XFILLER_38_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19645_ clknet_leaf_47_i_clk _00576_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16857_ _09462_ _09463_ vssd1 vssd1 vccd1 vccd1 _09464_ sky130_fd_sc_hd__nand2_1
XFILLER_66_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15808_ rbzero.traced_texa\[-9\] _08457_ _08459_ rbzero.wall_tracer.visualWallDist\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__a22o_1
X_16788_ _09354_ _09395_ vssd1 vssd1 vccd1 vccd1 _09396_ sky130_fd_sc_hd__xnor2_2
XFILLER_80_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19576_ clknet_leaf_30_i_clk _00507_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_15739_ _08321_ _08322_ _08420_ vssd1 vssd1 vccd1 vccd1 _08422_ sky130_fd_sc_hd__and3_1
X_18527_ _02481_ vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18458_ _02445_ vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__clkbuf_1
X_17409_ _01705_ _01706_ _01707_ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__o21ba_1
XFILLER_119_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20420_ net480 _01351_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20351_ net411 _01282_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20282_ net342 _01213_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[1\] sky130_fd_sc_hd__dfxtp_1
X_19035__209 clknet_1_1__leaf__02735_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__inv_2
XFILLER_161_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__02751_ clknet_0__02751_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02751_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11420_ _03652_ _04203_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__or2_1
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11351_ rbzero.debug_overlay.playerY\[-4\] _04089_ _04083_ rbzero.debug_overlay.playerY\[-7\]
+ _04135_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__a221o_1
XFILLER_192_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10302_ _03213_ vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14070_ rbzero.wall_tracer.trackDistX\[-5\] _06788_ _06798_ vssd1 vssd1 vccd1 vccd1
+ _00434_ sky130_fd_sc_hd__o21a_1
XFILLER_141_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11282_ gpout0.hpos\[5\] _04052_ _04054_ _04040_ vssd1 vssd1 vccd1 vccd1 _04067_
+ sky130_fd_sc_hd__or4b_2
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13021_ _05738_ _05736_ _05735_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__a21o_1
X_10233_ _03143_ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__clkbuf_4
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10164_ _03140_ vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10095_ _03104_ vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__clkbuf_1
X_14972_ _07653_ _07659_ vssd1 vssd1 vccd1 vccd1 _07660_ sky130_fd_sc_hd__xor2_1
X_17760_ _02018_ _02023_ _02026_ vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__nor3_1
XFILLER_48_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16711_ _09315_ _09316_ _09317_ vssd1 vssd1 vccd1 vccd1 _09319_ sky130_fd_sc_hd__and3_1
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13923_ _06615_ _06612_ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__or2_1
X_17691_ _01951_ _01963_ vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__nor2_1
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16642_ _08896_ _08889_ vssd1 vssd1 vccd1 vccd1 _09251_ sky130_fd_sc_hd__nor2_1
XFILLER_142_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19430_ _01919_ _01928_ _01927_ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13854_ _06559_ _06472_ vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12805_ _05354_ _05526_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__or2_1
X_16573_ _09181_ _09182_ vssd1 vssd1 vccd1 vccd1 _09183_ sky130_fd_sc_hd__nor2_1
XFILLER_16_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19361_ _02840_ _02841_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__and2b_1
X_13785_ _06504_ _06512_ _06529_ vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__and3_1
XFILLER_50_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10997_ gpout0.hpos\[2\] vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__clkinv_2
X_19140__304 clknet_1_1__leaf__02745_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__inv_2
X_15524_ _08204_ _08205_ _08207_ vssd1 vssd1 vccd1 vccd1 _08208_ sky130_fd_sc_hd__o21ai_1
X_18312_ _02390_ vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__clkbuf_1
XFILLER_187_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _05458_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__clkbuf_4
X_19292_ _02782_ _02783_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__xnor2_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ rbzero.spi_registers.new_vshift\[0\] _02348_ _02350_ _02314_ vssd1 vssd1
+ vccd1 vccd1 _00795_ sky130_fd_sc_hd__o211a_1
XFILLER_175_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15455_ _06771_ _06776_ _07893_ _06853_ vssd1 vssd1 vccd1 vccd1 _08140_ sky130_fd_sc_hd__a31o_1
XFILLER_176_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12667_ _05420_ _05422_ _05423_ _05333_ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__a31o_2
XFILLER_175_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14406_ _06966_ _07092_ vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__or2_1
XFILLER_198_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11618_ rbzero.tex_b1\[41\] rbzero.tex_b1\[40\] _03732_ vssd1 vssd1 vccd1 vccd1 _04399_
+ sky130_fd_sc_hd__mux2_1
X_18174_ rbzero.map_overlay.i_mapdy\[5\] _02291_ vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__or2_1
X_15386_ _08070_ vssd1 vssd1 vccd1 vccd1 _08071_ sky130_fd_sc_hd__clkbuf_4
XFILLER_168_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12598_ _05354_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__clkbuf_4
X_17125_ _09142_ _09231_ _09256_ _09229_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__or4_1
X_14337_ _06978_ _07024_ vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__or2_1
X_11549_ _03674_ _04326_ _04330_ _03704_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__a211o_1
XFILLER_117_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17056_ _08899_ _07961_ vssd1 vssd1 vccd1 vccd1 _09661_ sky130_fd_sc_hd__or2_1
X_14268_ rbzero.debug_overlay.playerY\[-4\] rbzero.debug_overlay.playerY\[-5\] _06922_
+ vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__or3_1
XFILLER_125_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16007_ _08619_ _08620_ vssd1 vssd1 vccd1 vccd1 _08621_ sky130_fd_sc_hd__nand2_1
Xclkbuf_0__02745_ _02745_ vssd1 vssd1 vccd1 vccd1 clknet_0__02745_ sky130_fd_sc_hd__clkbuf_16
X_13219_ _05925_ _05932_ _05975_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__a21oi_2
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _05075_ _05064_ _06885_ _06886_ vssd1 vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__a31o_2
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _02179_ vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16909_ _09423_ _09403_ _09514_ vssd1 vssd1 vccd1 vccd1 _09516_ sky130_fd_sc_hd__nand3_1
X_17889_ _02142_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__clkbuf_4
XFILLER_54_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19628_ clknet_leaf_45_i_clk _00559_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19559_ clknet_leaf_32_i_clk _00490_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20403_ net463 _01334_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20334_ net394 _01265_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20265_ net325 _01196_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20196_ net256 _01127_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10920_ rbzero.tex_r0\[25\] rbzero.tex_r0\[24\] _03690_ vssd1 vssd1 vccd1 vccd1 _03706_
+ sky130_fd_sc_hd__mux2_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19256__6 clknet_1_0__leaf__02433_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__inv_2
XFILLER_29_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02734_ clknet_0__02734_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02734_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_71_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18946__129 clknet_1_0__leaf__02726_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__inv_2
XFILLER_44_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10851_ rbzero.row_render.texu\[3\] rbzero.row_render.texu\[2\] rbzero.row_render.texu\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__nand3_1
XFILLER_71_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _06305_ _06326_ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__xor2_1
X_10782_ rbzero.traced_texVinit\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _03568_
+ sky130_fd_sc_hd__nand2_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _05198_ _05201_ _05257_ _05277_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__or4_2
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _07924_ _07926_ vssd1 vssd1 vccd1 vccd1 _07927_ sky130_fd_sc_hd__xor2_2
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ _05185_ _05208_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__nand2_4
XFILLER_123_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_61_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_200_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11403_ rbzero.tex_g0\[53\] rbzero.tex_g0\[52\] _03700_ vssd1 vssd1 vccd1 vccd1 _04187_
+ sky130_fd_sc_hd__mux2_1
XFILLER_184_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15171_ _07856_ _07857_ vssd1 vssd1 vccd1 vccd1 _07858_ sky130_fd_sc_hd__nor2_1
XFILLER_197_1140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12383_ _03479_ _04913_ _04914_ _05139_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__a31o_1
XFILLER_126_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14122_ rbzero.wall_tracer.stepDistX\[-2\] _06717_ _06825_ vssd1 vssd1 vccd1 vccd1
+ _06826_ sky130_fd_sc_hd__mux2_1
XFILLER_181_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11334_ rbzero.debug_overlay.facingX\[0\] _04079_ _04081_ rbzero.debug_overlay.facingX\[-9\]
+ _04118_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__a221o_1
XFILLER_181_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14053_ _05005_ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__clkbuf_4
XFILLER_158_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_76_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11265_ _04045_ _04049_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__xor2_1
XFILLER_107_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13004_ _05664_ _05684_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__xnor2_1
XFILLER_79_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10216_ _03168_ vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__clkbuf_1
X_18861_ _02693_ vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__clkbuf_1
X_11196_ rbzero.tex_r1\[26\] _03768_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__or2_1
XFILLER_122_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17812_ _08458_ _02066_ _02067_ _02076_ vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__a31o_1
XFILLER_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10147_ _03131_ vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__clkbuf_1
X_18792_ rbzero.debug_overlay.facingY\[-7\] _02645_ vssd1 vssd1 vccd1 vccd1 _02656_
+ sky130_fd_sc_hd__and2_1
X_14955_ _07541_ _07632_ _07637_ vssd1 vssd1 vccd1 vccd1 _07643_ sky130_fd_sc_hd__o21ai_1
X_17743_ _01985_ rbzero.wall_tracer.rayAddendX\[3\] vssd1 vssd1 vccd1 vccd1 _02012_
+ sky130_fd_sc_hd__and2_1
X_10078_ rbzero.tex_g1\[27\] rbzero.tex_g1\[28\] _03095_ vssd1 vssd1 vccd1 vccd1 _03096_
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13906_ _05325_ _06642_ vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__and2_1
X_17674_ rbzero.debug_overlay.vplaneX\[-7\] _01939_ vssd1 vssd1 vccd1 vccd1 _01949_
+ sky130_fd_sc_hd__nand2_1
XFILLER_78_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14886_ _07529_ _07570_ vssd1 vssd1 vccd1 vccd1 _07574_ sky130_fd_sc_hd__xor2_1
XFILLER_62_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19413_ _01707_ _01706_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__nor2_1
X_16625_ _09230_ _09232_ _09233_ vssd1 vssd1 vccd1 vccd1 _09234_ sky130_fd_sc_hd__o21ai_1
X_13837_ _06581_ _06584_ _06592_ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_14_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16556_ _07877_ _08803_ _09049_ vssd1 vssd1 vccd1 vccd1 _09166_ sky130_fd_sc_hd__o21ai_1
X_19344_ _02759_ _02826_ _02827_ _02319_ rbzero.texV\[2\] vssd1 vssd1 vccd1 vccd1
+ _01419_ sky130_fd_sc_hd__a32o_1
X_13768_ _06517_ _06523_ _06524_ vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__a21o_1
XFILLER_44_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15507_ rbzero.wall_tracer.visualWallDist\[9\] _07256_ vssd1 vssd1 vccd1 vccd1 _08191_
+ sky130_fd_sc_hd__nand2_4
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12719_ _05323_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__clkbuf_4
XFILLER_188_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16487_ _09095_ _09096_ vssd1 vssd1 vccd1 vccd1 _09097_ sky130_fd_sc_hd__nor2_1
XFILLER_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19275_ _02768_ _02769_ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__and2b_1
XFILLER_188_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13699_ _06408_ _06455_ vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__xor2_1
XFILLER_175_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15438_ _08120_ _08121_ vssd1 vssd1 vccd1 vccd1 _08123_ sky130_fd_sc_hd__or2_1
X_18226_ _03338_ _02338_ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_29_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_157_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18157_ rbzero.map_overlay.i_mapdx\[3\] _02292_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__or2_1
X_15369_ _08052_ _08053_ vssd1 vssd1 vccd1 vccd1 _08055_ sky130_fd_sc_hd__or2_1
XFILLER_157_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17108_ _09710_ _09711_ _09712_ vssd1 vssd1 vccd1 vccd1 _09713_ sky130_fd_sc_hd__a21oi_1
XFILLER_183_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18088_ rbzero.spi_registers.spi_cmd\[2\] rbzero.spi_registers.spi_cmd\[3\] _02245_
+ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__mux2_1
X_09930_ rbzero.tex_r0\[34\] rbzero.tex_r0\[33\] _03017_ vssd1 vssd1 vccd1 vccd1 _03018_
+ sky130_fd_sc_hd__mux2_1
X_17039_ _09021_ _09046_ vssd1 vssd1 vccd1 vccd1 _09644_ sky130_fd_sc_hd__nor2_1
XFILLER_171_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__02728_ _02728_ vssd1 vssd1 vccd1 vccd1 clknet_0__02728_ sky130_fd_sc_hd__clkbuf_16
X_20050_ clknet_leaf_82_i_clk _00981_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[66\]
+ sky130_fd_sc_hd__dfxtp_1
X_09861_ rbzero.tex_r1\[0\] rbzero.tex_r1\[1\] _02976_ vssd1 vssd1 vccd1 vccd1 _02980_
+ sky130_fd_sc_hd__mux2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09792_ rbzero.tex_r1\[33\] rbzero.tex_r1\[34\] _02943_ vssd1 vssd1 vccd1 vccd1 _02944_
+ sky130_fd_sc_hd__mux2_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20317_ net377 _01248_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11050_ gpout0.vpos\[6\] _03347_ rbzero.debug_overlay.playerX\[0\] _03462_ _03835_
+ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__o221a_1
X_20248_ net308 _01179_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10001_ rbzero.tex_g1\[63\] net48 _02976_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__mux2_1
XFILLER_88_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20179_ net239 _01110_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19013__189 clknet_1_1__leaf__02733_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__inv_2
XFILLER_76_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14740_ _07396_ _07398_ vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__xnor2_1
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ _04724_ _04725_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__and2_1
XFILLER_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_106 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_106/HI zeros[15]
+ sky130_fd_sc_hd__conb_1
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_117 vssd1 vssd1 vccd1 vccd1 ones[10] top_ew_algofoogle_117/LO sky130_fd_sc_hd__conb_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10903_ _03669_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__buf_6
XFILLER_72_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ _07341_ _07358_ vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__nand2_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ _03910_ _04622_ _04625_ net69 vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__a22o_1
XFILLER_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16410_ _08108_ vssd1 vssd1 vccd1 vccd1 _09021_ sky130_fd_sc_hd__clkbuf_4
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13622_ _06358_ _06377_ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__nor2_1
X_10834_ _03556_ _03613_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__and2_2
X_17390_ _03369_ _01691_ _08506_ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__mux2_1
XFILLER_77_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16341_ _08826_ _08827_ _08829_ vssd1 vssd1 vccd1 vccd1 _08953_ sky130_fd_sc_hd__o21a_2
XFILLER_13_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13553_ _06259_ _06264_ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10765_ _03548_ _03547_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__nand2_1
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12504_ _05118_ _05239_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__xor2_2
XFILLER_185_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16272_ _08787_ _08796_ vssd1 vssd1 vccd1 vccd1 _08884_ sky130_fd_sc_hd__nand2_1
XFILLER_73_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13484_ _06103_ _05988_ _06239_ _06240_ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__o31ai_2
XFILLER_200_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10696_ _03482_ _03486_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__nor2_1
XFILLER_185_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15223_ _07886_ _07909_ vssd1 vssd1 vccd1 vccd1 _07910_ sky130_fd_sc_hd__xnor2_2
X_18011_ rbzero.pov.spi_buffer\[58\] rbzero.pov.ready_buffer\[58\] _02197_ vssd1 vssd1
+ vccd1 vccd1 _02207_ sky130_fd_sc_hd__mux2_1
X_12435_ _05190_ _05191_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__xnor2_2
XFILLER_139_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15154_ _07838_ _07840_ vssd1 vssd1 vccd1 vccd1 _07841_ sky130_fd_sc_hd__xor2_1
X_12366_ _05122_ _05038_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__nor2_1
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14105_ rbzero.wall_tracer.stepDistX\[-10\] _06649_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _06817_ sky130_fd_sc_hd__mux2_1
X_11317_ rbzero.debug_overlay.vplaneX\[-4\] vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__clkbuf_4
XFILLER_180_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19962_ net191 _00893_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[42\] sky130_fd_sc_hd__dfxtp_1
X_15085_ _07771_ _07772_ vssd1 vssd1 vccd1 vccd1 _07773_ sky130_fd_sc_hd__nor2_1
XFILLER_4_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12297_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] _05053_
+ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__o21a_1
X_14036_ _06097_ _05305_ vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__nor2_2
XFILLER_141_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11248_ _03500_ _04032_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__nor2_1
XFILLER_171_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19893_ clknet_leaf_18_i_clk _00824_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_110_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18844_ rbzero.pov.ready_buffer\[3\] _02666_ _02684_ _02675_ vssd1 vssd1 vccd1 vccd1
+ _01062_ sky130_fd_sc_hd__a211o_1
XFILLER_45_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11179_ rbzero.tex_r1\[3\] _03936_ _03963_ _03726_ vssd1 vssd1 vccd1 vccd1 _03964_
+ sky130_fd_sc_hd__o211a_1
XFILLER_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18775_ rbzero.debug_overlay.facingX\[-4\] _02645_ vssd1 vssd1 vccd1 vccd1 _02647_
+ sky130_fd_sc_hd__and2_1
X_15987_ _08352_ _08599_ _08600_ vssd1 vssd1 vccd1 vccd1 _08601_ sky130_fd_sc_hd__a21oi_1
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17726_ _01996_ vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__inv_2
X_14938_ _07623_ _07624_ _07625_ vssd1 vssd1 vccd1 vccd1 _07626_ sky130_fd_sc_hd__o21a_1
XFILLER_36_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17657_ _04102_ rbzero.wall_tracer.rayAddendX\[-4\] vssd1 vssd1 vccd1 vccd1 _01933_
+ sky130_fd_sc_hd__or2_1
X_14869_ _07554_ _07556_ vssd1 vssd1 vccd1 vccd1 _07557_ sky130_fd_sc_hd__or2b_1
XFILLER_51_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16608_ _09216_ vssd1 vssd1 vccd1 vccd1 _09217_ sky130_fd_sc_hd__inv_2
XFILLER_51_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17588_ _01871_ _01859_ _01873_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19327_ _02806_ _02810_ _02811_ _02812_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__o211a_1
X_16539_ _09138_ _09148_ vssd1 vssd1 vccd1 vccd1 _09149_ sky130_fd_sc_hd__xnor2_1
XFILLER_177_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19258_ gpout5.clk_div\[1\] gpout5.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__nand2_1
XFILLER_31_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18209_ _03338_ _02326_ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__or2_1
XFILLER_191_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09913_ rbzero.tex_r0\[42\] rbzero.tex_r0\[41\] _03006_ vssd1 vssd1 vccd1 vccd1 _03009_
+ sky130_fd_sc_hd__mux2_1
X_20102_ clknet_leaf_90_i_clk _01033_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_132_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20033_ clknet_leaf_86_i_clk _00964_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09844_ rbzero.tex_r1\[8\] rbzero.tex_r1\[9\] _02965_ vssd1 vssd1 vccd1 vccd1 _02971_
+ sky130_fd_sc_hd__mux2_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09775_ rbzero.tex_r1\[41\] rbzero.tex_r1\[42\] _02932_ vssd1 vssd1 vccd1 vccd1 _02935_
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__02433_ clknet_0__02433_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02433_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19201__359 clknet_1_0__leaf__02751_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__inv_2
XFILLER_195_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10550_ _03345_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__inv_2
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10481_ rbzero.tex_b0\[28\] rbzero.tex_b0\[27\] _03302_ vssd1 vssd1 vccd1 vccd1 _03307_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12220_ _04972_ rbzero.wall_tracer.trackDistX\[-6\] rbzero.wall_tracer.trackDistX\[-7\]
+ _04973_ _04981_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__a221o_1
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12151_ _04870_ _04873_ _04912_ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__o21bai_1
XFILLER_155_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11102_ rbzero.debug_overlay.playerX\[-3\] gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1
+ _03888_ sky130_fd_sc_hd__xnor2_1
XFILLER_150_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12082_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] vssd1
+ vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__or2_1
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11033_ _02903_ _03793_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__nor2_1
X_15910_ _08524_ _07815_ vssd1 vssd1 vccd1 vccd1 _08532_ sky130_fd_sc_hd__and2_1
X_16890_ _09478_ _09479_ _09495_ vssd1 vssd1 vccd1 vccd1 _09497_ sky130_fd_sc_hd__nand3_1
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ _08469_ _08470_ vssd1 vssd1 vccd1 vccd1 _08471_ sky130_fd_sc_hd__nor2_1
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18560_ _02498_ vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ _05484_ _05473_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__nand2_1
X_15772_ _08445_ vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__clkbuf_1
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17511_ _01799_ _01800_ _01797_ _01798_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__o211ai_1
X_14723_ _06872_ _07273_ _07410_ vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__nor3_1
X_11935_ _04532_ _04709_ _04680_ net48 vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__a31o_1
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18491_ _02462_ vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17442_ _01726_ _01729_ _01737_ vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__o21ai_1
XFILLER_45_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14654_ _07301_ _07305_ vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__xnor2_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11866_ net50 _04622_ _04641_ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__a21o_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _06289_ _06338_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__xnor2_1
X_10817_ _03570_ _03601_ _03602_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__o21a_4
X_14585_ _07037_ vssd1 vssd1 vccd1 vccd1 _07273_ sky130_fd_sc_hd__buf_4
X_17373_ rbzero.spi_registers.new_mapd\[15\] rbzero.spi_registers.spi_buffer\[15\]
+ _01662_ vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__mux2_1
X_11797_ _03910_ _04566_ _04568_ net69 _04573_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__a221o_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16324_ _08932_ _08934_ vssd1 vssd1 vccd1 vccd1 _08936_ sky130_fd_sc_hd__and2_1
X_13536_ _06103_ _05992_ _06291_ _06292_ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__o31ai_2
XFILLER_186_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10748_ _03530_ _03532_ _03533_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__nor3_2
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16255_ _07993_ _07333_ _07787_ _08643_ vssd1 vssd1 vccd1 vccd1 _08867_ sky130_fd_sc_hd__o22ai_1
X_19043_ clknet_1_0__leaf__02732_ vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__buf_1
XFILLER_174_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13467_ _06208_ _06222_ _06223_ vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__and3_1
XFILLER_199_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10679_ _03473_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__buf_4
X_15206_ _06759_ _06764_ _06767_ _07165_ vssd1 vssd1 vccd1 vccd1 _07893_ sky130_fd_sc_hd__nor4_4
X_12418_ _05167_ _05168_ _05174_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__o21ba_1
XFILLER_161_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16186_ _07661_ _08678_ vssd1 vssd1 vccd1 vccd1 _08799_ sky130_fd_sc_hd__or2_1
X_13398_ _05902_ _05903_ vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__xnor2_1
XFILLER_182_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15137_ _06914_ vssd1 vssd1 vccd1 vccd1 _07825_ sky130_fd_sc_hd__clkbuf_4
XFILLER_99_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12349_ _05041_ _05042_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__and2b_1
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19945_ net174 _00876_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15068_ _04841_ rbzero.wall_tracer.stepDistX\[4\] _07171_ _07172_ vssd1 vssd1 vccd1
+ vccd1 _07756_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_99_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14019_ _06760_ vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19876_ clknet_leaf_18_i_clk _00807_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18827_ rbzero.debug_overlay.vplaneX\[-3\] _02660_ vssd1 vssd1 vccd1 vccd1 _02676_
+ sky130_fd_sc_hd__or2_1
XFILLER_56_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18758_ _02634_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__buf_2
XFILLER_67_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17709_ _04100_ rbzero.debug_overlay.vplaneX\[-9\] _01980_ vssd1 vssd1 vccd1 vccd1
+ _01981_ sky130_fd_sc_hd__a21oi_1
XFILLER_64_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18689_ net40 _02532_ _02262_ vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09827_ rbzero.tex_r1\[16\] rbzero.tex_r1\[17\] _02954_ vssd1 vssd1 vccd1 vccd1 _02962_
+ sky130_fd_sc_hd__mux2_1
X_20016_ clknet_leaf_92_i_clk _00947_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09758_ rbzero.tex_r1\[49\] rbzero.tex_r1\[50\] _02921_ vssd1 vssd1 vccd1 vccd1 _02926_
+ sky130_fd_sc_hd__mux2_1
XFILLER_100_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11720_ _04489_ _04492_ _04497_ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__and3_1
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _04423_ _04431_ _03685_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__a21o_1
XFILLER_42_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10602_ _03395_ _03343_ _03396_ _03397_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__a31o_1
X_14370_ _07056_ _07057_ vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__nor2_1
X_11582_ _04361_ _04362_ _04363_ _04192_ _03607_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__o221a_1
XFILLER_11_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13321_ _06076_ _06077_ vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__nand2_1
X_10533_ rbzero.tex_b0\[3\] rbzero.tex_b0\[2\] _03324_ vssd1 vssd1 vccd1 vccd1 _03334_
+ sky130_fd_sc_hd__mux2_1
XFILLER_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16040_ _08651_ _08652_ vssd1 vssd1 vccd1 vccd1 _08654_ sky130_fd_sc_hd__and2_1
XFILLER_127_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13252_ _05355_ _06008_ _05593_ _05301_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__o22a_1
X_10464_ rbzero.tex_b0\[36\] rbzero.tex_b0\[35\] _03291_ vssd1 vssd1 vccd1 vccd1 _03298_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12203_ _04963_ rbzero.wall_tracer.trackDistX\[0\] _04964_ rbzero.wall_tracer.trackDistX\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__a22o_1
XFILLER_109_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13183_ _05938_ _05910_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__or2b_1
X_10395_ rbzero.tex_b1\[4\] rbzero.tex_b1\[5\] _03254_ vssd1 vssd1 vccd1 vccd1 _03262_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12134_ _04859_ _04895_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__nand2_1
XFILLER_151_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19019__195 clknet_1_0__leaf__02733_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__inv_2
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17991_ _02196_ vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19730_ clknet_leaf_94_i_clk _00661_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16942_ _09046_ _09547_ vssd1 vssd1 vccd1 vccd1 _09548_ sky130_fd_sc_hd__nor2_1
X_12065_ _04833_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__buf_4
XFILLER_81_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11016_ rbzero.row_render.size\[4\] _03773_ rbzero.row_render.size\[5\] vssd1 vssd1
+ vccd1 vccd1 _03802_ sky130_fd_sc_hd__o21ai_1
X_19661_ clknet_leaf_4_i_clk _00592_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_16873_ _09009_ _09007_ _09256_ _09039_ vssd1 vssd1 vccd1 vccd1 _09480_ sky130_fd_sc_hd__nor4_1
XFILLER_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18612_ _02525_ vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15824_ rbzero.traced_texa\[4\] _08461_ _08462_ rbzero.wall_tracer.visualWallDist\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__a22o_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19592_ clknet_leaf_40_i_clk _00523_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18543_ rbzero.pov.spi_buffer\[40\] rbzero.pov.spi_buffer\[41\] _02488_ vssd1 vssd1
+ vccd1 vccd1 _02490_ sky130_fd_sc_hd__mux2_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ _05680_ _05723_ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__xor2_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15755_ _03337_ _03506_ vssd1 vssd1 vccd1 vccd1 _08437_ sky130_fd_sc_hd__or2_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14706_ _06949_ _07005_ vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__or2_1
X_11918_ _04670_ _04692_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__nand2_1
X_18474_ _02453_ vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15686_ _08367_ _08368_ vssd1 vssd1 vccd1 vccd1 _08369_ sky130_fd_sc_hd__nand2_1
X_12898_ _05516_ _05474_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__nor2_1
XFILLER_33_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__or2_1
XFILLER_21_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14637_ _07323_ _07324_ vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__nand2_1
X_11849_ net10 net9 vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__and2b_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14568_ _06855_ vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__clkbuf_8
X_17356_ _01670_ vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16307_ _08917_ _08918_ vssd1 vssd1 vccd1 vccd1 _08919_ sky130_fd_sc_hd__and2_1
X_13519_ _06273_ _06275_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__or2b_1
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17287_ rbzero.wall_tracer.trackDistY\[3\] _01558_ _01615_ _09081_ vssd1 vssd1 vccd1
+ vccd1 _00574_ sky130_fd_sc_hd__o22a_1
X_14499_ _07182_ _07184_ _07186_ vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__a21boi_1
X_16238_ _07984_ _07865_ _07959_ _08070_ vssd1 vssd1 vccd1 vccd1 _08850_ sky130_fd_sc_hd__or4_1
XFILLER_134_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16169_ _08772_ _08781_ vssd1 vssd1 vccd1 vccd1 _08782_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19928_ net157 _00859_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_130_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19859_ clknet_leaf_21_i_clk _00790_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19234__9 clknet_1_1__leaf__02754_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__inv_2
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20496_ clknet_leaf_44_i_clk _01427_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10180_ _03149_ vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13870_ _05271_ _06626_ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__nor2_1
XFILLER_46_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12821_ _05355_ _05551_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__nor2_1
XFILLER_74_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15540_ _06875_ _07735_ vssd1 vssd1 vccd1 vccd1 _08224_ sky130_fd_sc_hd__nor2_1
X_19207__365 clknet_1_1__leaf__02751_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__inv_2
X_12752_ _05507_ _05508_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11703_ _03505_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__inv_2
X_15471_ _08154_ _08155_ vssd1 vssd1 vccd1 vccd1 _08156_ sky130_fd_sc_hd__nor2_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _05336_ _05337_ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__nand2_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _07101_ _07109_ vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__or2_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _01541_ _01543_ _01542_ vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__a21boi_1
X_11634_ _03679_ _04402_ _04406_ _04410_ _04414_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__o32a_1
XFILLER_30_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18190_ rbzero.spi_registers.new_leak\[1\] _02310_ _02313_ _02314_ vssd1 vssd1 vccd1
+ vccd1 _00778_ sky130_fd_sc_hd__o211a_1
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17141_ _09662_ _01484_ vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__xnor2_2
X_14353_ _07006_ _07039_ _07040_ vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__or3_1
X_11565_ _04179_ _04342_ _04346_ _03624_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__a211o_1
XFILLER_195_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13304_ _06035_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__clkbuf_4
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17072_ rbzero.wall_tracer.visualWallDist\[4\] _07256_ _07173_ _09675_ _09676_ vssd1
+ vssd1 vccd1 vccd1 _09677_ sky130_fd_sc_hd__a41o_1
X_10516_ _03325_ vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__02730_ clknet_0__02730_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02730_
+ sky130_fd_sc_hd__clkbuf_16
X_14284_ _06967_ _06971_ vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__nand2_1
X_11496_ _04277_ _04278_ _03917_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__mux2_1
XFILLER_183_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16023_ _08370_ _08371_ _08373_ vssd1 vssd1 vccd1 vccd1 _08637_ sky130_fd_sc_hd__o21ai_1
X_13235_ _05991_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__clkbuf_4
X_10447_ rbzero.tex_b0\[44\] rbzero.tex_b0\[43\] _03280_ vssd1 vssd1 vccd1 vccd1 _03289_
+ sky130_fd_sc_hd__mux2_1
XFILLER_109_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13166_ _05921_ _05922_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__nand2_1
X_10378_ rbzero.tex_b1\[12\] rbzero.tex_b1\[13\] _03243_ vssd1 vssd1 vccd1 vccd1 _03253_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12117_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[10\] vssd1
+ vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__nor2_1
X_17974_ rbzero.pov.spi_buffer\[40\] rbzero.pov.ready_buffer\[40\] _02186_ vssd1 vssd1
+ vccd1 vccd1 _02188_ sky130_fd_sc_hd__mux2_1
X_13097_ _05760_ _05765_ _05853_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__a21o_1
X_19713_ clknet_leaf_2_i_clk _00644_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16925_ _09529_ _09530_ vssd1 vssd1 vccd1 vccd1 _09531_ sky130_fd_sc_hd__nor2_1
X_12048_ net34 net33 gpout5.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__and3_1
XFILLER_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19644_ clknet_leaf_48_i_clk _00575_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16856_ _09461_ _09460_ vssd1 vssd1 vccd1 vccd1 _09463_ sky130_fd_sc_hd__or2b_1
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15807_ _08458_ vssd1 vssd1 vccd1 vccd1 _08459_ sky130_fd_sc_hd__buf_2
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19575_ clknet_leaf_30_i_clk _00506_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_16787_ _09393_ _09394_ vssd1 vssd1 vccd1 vccd1 _09395_ sky130_fd_sc_hd__xor2_2
XFILLER_81_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13999_ _06742_ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__clkinv_2
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18526_ rbzero.pov.spi_buffer\[32\] rbzero.pov.spi_buffer\[33\] _02477_ vssd1 vssd1
+ vccd1 vccd1 _02481_ sky130_fd_sc_hd__mux2_1
X_15738_ _08321_ _08322_ _08420_ vssd1 vssd1 vccd1 vccd1 _08421_ sky130_fd_sc_hd__a21oi_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18457_ rbzero.pov.mosi rbzero.pov.spi_buffer\[0\] _02444_ vssd1 vssd1 vccd1 vccd1
+ _02445_ sky130_fd_sc_hd__mux2_1
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15669_ _08240_ _08324_ _08351_ vssd1 vssd1 vccd1 vccd1 _08352_ sky130_fd_sc_hd__a21o_1
XFILLER_34_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17408_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.wall_tracer.rayAddendY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__and2_1
XFILLER_92_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17339_ _01659_ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__inv_2
XFILLER_140_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20350_ net410 _01281_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19009_ clknet_1_1__leaf__04486_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__buf_1
XFILLER_106_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20281_ net341 _01212_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__02750_ clknet_0__02750_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02750_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_56_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18433__73 clknet_1_0__leaf__02438_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__inv_2
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11350_ rbzero.debug_overlay.playerY\[5\] _04125_ _03519_ _03854_ vssd1 vssd1 vccd1
+ vccd1 _04135_ sky130_fd_sc_hd__a211o_1
XFILLER_138_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10301_ rbzero.tex_b1\[49\] rbzero.tex_b1\[50\] _03210_ vssd1 vssd1 vccd1 vccd1 _03213_
+ sky130_fd_sc_hd__mux2_1
XFILLER_180_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11281_ _04051_ _04065_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__nor2_1
XFILLER_106_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20479_ clknet_leaf_63_i_clk _01410_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13020_ _05738_ _05735_ _05736_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__nand3_1
XFILLER_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10232_ _03176_ vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10163_ rbzero.tex_g0\[51\] rbzero.tex_g0\[50\] _03132_ vssd1 vssd1 vccd1 vccd1 _03140_
+ sky130_fd_sc_hd__mux2_1
XFILLER_121_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10094_ rbzero.tex_g1\[19\] rbzero.tex_g1\[20\] _03095_ vssd1 vssd1 vccd1 vccd1 _03104_
+ sky130_fd_sc_hd__mux2_1
X_14971_ _07654_ _07658_ _07656_ vssd1 vssd1 vccd1 vccd1 _07659_ sky130_fd_sc_hd__a21oi_1
XFILLER_59_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16710_ _09315_ _09316_ _09317_ vssd1 vssd1 vccd1 vccd1 _09318_ sky130_fd_sc_hd__a21oi_2
X_13922_ _05310_ vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__buf_2
X_17690_ _01952_ _01954_ vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__nor2_1
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16641_ _09248_ _09249_ vssd1 vssd1 vccd1 vccd1 _09250_ sky130_fd_sc_hd__nand2_1
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13853_ _06601_ _06609_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__and2_1
XFILLER_16_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19360_ rbzero.traced_texa\[5\] rbzero.texV\[5\] vssd1 vssd1 vccd1 vccd1 _02841_
+ sky130_fd_sc_hd__nand2_1
X_12804_ _05491_ _05560_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__and2_1
X_16572_ _09005_ _09064_ _09063_ vssd1 vssd1 vccd1 vccd1 _09182_ sky130_fd_sc_hd__a21oi_1
XFILLER_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13784_ _06539_ _06540_ vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__or2_1
X_10996_ _03781_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__buf_4
XFILLER_43_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18311_ rbzero.spi_registers.new_other\[1\] rbzero.spi_registers.spi_buffer\[1\]
+ _02388_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__mux2_1
X_15523_ _08078_ _08206_ vssd1 vssd1 vccd1 vccd1 _08207_ sky130_fd_sc_hd__nand2_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _05488_ _05489_ _05490_ _05491_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__o31a_2
XFILLER_15_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19291_ _02777_ _02779_ _02778_ vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__o21bai_1
XFILLER_188_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18923__108 clknet_1_0__leaf__02724_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__inv_2
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ rbzero.spi_registers.vshift\[0\] _02349_ vssd1 vssd1 vccd1 vccd1 _02350_
+ sky130_fd_sc_hd__or2_1
XFILLER_187_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12666_ _05261_ _05349_ _05371_ _05395_ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__o211ai_1
X_15454_ _06771_ _07893_ _06777_ vssd1 vssd1 vccd1 vccd1 _08139_ sky130_fd_sc_hd__a21boi_1
XFILLER_187_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11617_ _03621_ _04397_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__nor2_1
X_14405_ _06968_ _07092_ vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__nor2_1
XFILLER_129_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18173_ rbzero.spi_registers.new_mapd\[8\] _02289_ _02304_ _02301_ vssd1 vssd1 vccd1
+ vccd1 _00771_ sky130_fd_sc_hd__o211a_1
X_15385_ _08069_ vssd1 vssd1 vccd1 vccd1 _08070_ sky130_fd_sc_hd__buf_2
XFILLER_156_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12597_ _05328_ _05353_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__nor2_1
XFILLER_184_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17124_ _08888_ _08317_ _09670_ _09668_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__a31o_1
XFILLER_190_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11548_ _04192_ _04327_ _04328_ _04329_ _04179_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__o221a_1
X_14336_ _07019_ _07020_ _07023_ _04948_ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__a22o_4
XFILLER_144_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17055_ _09539_ _09558_ _09659_ vssd1 vssd1 vccd1 vccd1 _09660_ sky130_fd_sc_hd__a21bo_1
XFILLER_144_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14267_ _06949_ _06954_ vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__or2_1
X_11479_ rbzero.tex_g1\[8\] _03618_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__and2_1
Xclkbuf_0__02744_ _02744_ vssd1 vssd1 vccd1 vccd1 clknet_0__02744_ sky130_fd_sc_hd__clkbuf_16
X_16006_ _07084_ _07787_ _08339_ vssd1 vssd1 vccd1 vccd1 _08620_ sky130_fd_sc_hd__o21ai_1
X_13218_ _05882_ _05933_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__and2b_1
XFILLER_83_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14198_ _05062_ _05060_ _05061_ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__a21oi_1
XFILLER_87_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _05900_ _05905_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__nand2_1
XFILLER_48_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ rbzero.pov.spi_buffer\[32\] rbzero.pov.ready_buffer\[32\] _02175_ vssd1 vssd1
+ vccd1 vccd1 _02179_ sky130_fd_sc_hd__mux2_1
XFILLER_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16908_ _09423_ _09403_ _09514_ vssd1 vssd1 vccd1 vccd1 _09515_ sky130_fd_sc_hd__a21oi_1
XFILLER_66_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17888_ _02141_ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__clkbuf_4
XFILLER_66_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19627_ clknet_leaf_45_i_clk _00558_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_16839_ _07766_ _08130_ _09231_ _09229_ vssd1 vssd1 vccd1 vccd1 _09446_ sky130_fd_sc_hd__or4_1
XFILLER_66_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19558_ clknet_leaf_12_i_clk _00489_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_94_1120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18509_ rbzero.pov.spi_buffer\[24\] rbzero.pov.spi_buffer\[25\] _02466_ vssd1 vssd1
+ vccd1 vccd1 _02472_ sky130_fd_sc_hd__mux2_1
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19489_ clknet_leaf_61_i_clk _00435_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20402_ net462 _01333_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20333_ net393 _01264_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20264_ net324 _01195_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20195_ net255 _01126_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_130_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02733_ clknet_0__02733_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02733_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ _03627_ _03634_ _03635_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__or3_1
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10781_ _03550_ _03558_ _03566_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__o21a_1
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12520_ _05221_ _05222_ _05223_ _05254_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__or4_1
XFILLER_201_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _05198_ _05201_ _05207_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__and3b_1
XFILLER_200_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11402_ _03688_ _04160_ _04168_ _04185_ _03719_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__a311o_1
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15170_ _07270_ vssd1 vssd1 vccd1 vccd1 _07857_ sky130_fd_sc_hd__clkbuf_4
X_12382_ rbzero.wall_tracer.visualWallDist\[0\] _05067_ _03488_ vssd1 vssd1 vccd1
+ vccd1 _05139_ sky130_fd_sc_hd__a21o_1
XFILLER_181_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14121_ _04833_ vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__buf_4
XFILLER_126_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11333_ rbzero.debug_overlay.facingX\[-7\] _04083_ _04085_ rbzero.debug_overlay.facingX\[-5\]
+ _04117_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__a221o_1
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14052_ rbzero.wall_tracer.visualWallDist\[-11\] vssd1 vssd1 vccd1 vccd1 _06787_
+ sky130_fd_sc_hd__buf_4
XFILLER_107_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11264_ gpout0.hpos\[8\] _04048_ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13003_ _05726_ _05759_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__nor2_1
X_10215_ rbzero.tex_g0\[27\] rbzero.tex_g0\[26\] _03166_ vssd1 vssd1 vccd1 vccd1 _03168_
+ sky130_fd_sc_hd__mux2_1
X_18860_ _02143_ _02692_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__and2_1
X_11195_ rbzero.tex_r1\[28\] _03661_ _03936_ _03979_ vssd1 vssd1 vccd1 vccd1 _03980_
+ sky130_fd_sc_hd__a31o_1
XFILLER_122_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17811_ _03340_ _02074_ _02075_ _08448_ rbzero.wall_tracer.rayAddendX\[7\] vssd1
+ vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__a32o_1
X_10146_ rbzero.tex_g0\[59\] rbzero.tex_g0\[58\] _03050_ vssd1 vssd1 vccd1 vccd1 _03131_
+ sky130_fd_sc_hd__mux2_1
XFILLER_121_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18791_ rbzero.pov.ready_buffer\[23\] _02636_ _02655_ _02643_ vssd1 vssd1 vccd1 vccd1
+ _01038_ sky130_fd_sc_hd__o211a_1
XFILLER_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17742_ _01985_ rbzero.wall_tracer.rayAddendX\[2\] _01990_ vssd1 vssd1 vccd1 vccd1
+ _02011_ sky130_fd_sc_hd__o21bai_1
XFILLER_94_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10077_ _03072_ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__clkbuf_4
X_14954_ _07611_ _07641_ vssd1 vssd1 vccd1 vccd1 _07642_ sky130_fd_sc_hd__xor2_1
XFILLER_134_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13905_ _06659_ vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__clkbuf_1
X_17673_ rbzero.debug_overlay.vplaneX\[-7\] _01939_ vssd1 vssd1 vccd1 vccd1 _01948_
+ sky130_fd_sc_hd__or2_1
X_14885_ _07571_ _07572_ vssd1 vssd1 vccd1 vccd1 _07573_ sky130_fd_sc_hd__and2b_1
X_19412_ rbzero.wall_tracer.rayAddendY\[-9\] _08449_ _02873_ vssd1 vssd1 vccd1 vccd1
+ _01441_ sky130_fd_sc_hd__a21o_1
X_16624_ _07878_ _08252_ _09231_ _09229_ vssd1 vssd1 vccd1 vccd1 _09233_ sky130_fd_sc_hd__or4_1
XFILLER_165_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19064__236 clknet_1_0__leaf__02737_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__inv_2
X_13836_ _06581_ _06592_ vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__xor2_2
X_18412__54 clknet_1_1__leaf__02436_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__inv_2
XFILLER_51_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19343_ _02822_ _02823_ _02824_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__a21o_1
X_16555_ _08807_ _09052_ vssd1 vssd1 vccd1 vccd1 _09165_ sky130_fd_sc_hd__nand2_1
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10979_ _03686_ _03720_ _03746_ _03763_ _03764_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__o221a_1
X_13767_ _06518_ _06522_ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__and2b_1
XFILLER_189_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15506_ _08096_ _08113_ _08189_ vssd1 vssd1 vccd1 vccd1 _08190_ sky130_fd_sc_hd__a21bo_1
XFILLER_189_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12718_ _05473_ _05474_ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__nor2_1
X_19274_ rbzero.traced_texa\[-9\] rbzero.texV\[-9\] vssd1 vssd1 vccd1 vccd1 _02769_
+ sky130_fd_sc_hd__nand2_1
X_16486_ _09002_ _09093_ _09094_ vssd1 vssd1 vccd1 vccd1 _09096_ sky130_fd_sc_hd__and3_1
XFILLER_148_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13698_ _06121_ _06070_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__nor2_1
XFILLER_188_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18225_ rbzero.color_floor\[1\] rbzero.spi_registers.new_floor\[1\] _02335_ vssd1
+ vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__mux2_1
X_15437_ _08120_ _08121_ vssd1 vssd1 vccd1 vccd1 _08122_ sky130_fd_sc_hd__nand2_1
XFILLER_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12649_ _05219_ _05305_ _05302_ _05306_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__or4_1
XFILLER_175_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18156_ rbzero.spi_registers.new_mapd\[12\] _02290_ _02295_ _02275_ vssd1 vssd1 vccd1
+ vccd1 _00763_ sky130_fd_sc_hd__o211a_1
X_15368_ _08052_ _08053_ vssd1 vssd1 vccd1 vccd1 _08054_ sky130_fd_sc_hd__nand2_1
XFILLER_190_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17107_ _09623_ _09625_ _09624_ vssd1 vssd1 vccd1 vccd1 _09712_ sky130_fd_sc_hd__a21bo_1
X_14319_ _07006_ vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__clkbuf_4
XFILLER_183_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18087_ _02248_ vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__clkbuf_1
X_15299_ _07984_ _07281_ _07862_ _07861_ vssd1 vssd1 vccd1 vccd1 _07985_ sky130_fd_sc_hd__o31a_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17038_ _09547_ _09642_ vssd1 vssd1 vccd1 vccd1 _09643_ sky130_fd_sc_hd__nand2_1
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__02727_ _02727_ vssd1 vssd1 vccd1 vccd1 clknet_0__02727_ sky130_fd_sc_hd__clkbuf_16
X_09860_ _02979_ vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _02909_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__clkbuf_4
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20316_ net376 _01247_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20247_ net307 _01178_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10000_ _03054_ vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20178_ net238 _01109_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_130_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09989_ _03048_ vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11951_ net30 net29 vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__nor2_2
XFILLER_85_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xtop_ew_algofoogle_107 vssd1 vssd1 vccd1 vccd1 ones[0] top_ew_algofoogle_107/LO sky130_fd_sc_hd__conb_1
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10902_ _03687_ vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__buf_6
XFILLER_45_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_118 vssd1 vssd1 vccd1 vccd1 ones[11] top_ew_algofoogle_118/LO sky130_fd_sc_hd__conb_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14670_ _07355_ _07356_ _07357_ vssd1 vssd1 vccd1 vccd1 _07358_ sky130_fd_sc_hd__a21oi_1
X_11882_ _04645_ _04651_ _04655_ _04657_ net13 vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__o221a_1
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10833_ rbzero.row_render.texu\[0\] _03607_ _03612_ _03618_ _03538_ vssd1 vssd1 vccd1
+ vccd1 _03619_ sky130_fd_sc_hd__a41o_1
X_13621_ _06358_ _06377_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__xor2_1
XFILLER_26_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16340_ _08725_ _08951_ vssd1 vssd1 vccd1 vccd1 _08952_ sky130_fd_sc_hd__xnor2_4
XFILLER_73_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10764_ _03546_ _03549_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__nor2_1
X_13552_ _06295_ _06301_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__xor2_1
XFILLER_34_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12503_ _05256_ _05198_ _05257_ _05259_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__or4_1
XFILLER_186_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16271_ _08772_ _08781_ _08779_ vssd1 vssd1 vccd1 vccd1 _08883_ sky130_fd_sc_hd__a21o_1
X_13483_ _05862_ _06061_ _06238_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__or3_1
XFILLER_9_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10695_ _03340_ vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__buf_4
XFILLER_201_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18010_ _02206_ vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__clkbuf_1
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15222_ _07906_ _07908_ vssd1 vssd1 vccd1 vccd1 _07909_ sky130_fd_sc_hd__xor2_2
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12434_ _05133_ _05146_ _05187_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__o21ai_1
XFILLER_201_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15153_ _06866_ _07839_ vssd1 vssd1 vccd1 vccd1 _07840_ sky130_fd_sc_hd__nor2_1
X_12365_ rbzero.debug_overlay.facingX\[-7\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__and2_1
XFILLER_154_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11316_ rbzero.debug_overlay.vplaneX\[-8\] _04090_ _04085_ _04100_ vssd1 vssd1 vccd1
+ vccd1 _04101_ sky130_fd_sc_hd__a22o_1
X_14104_ _06816_ vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19961_ net190 _00892_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[41\] sky130_fd_sc_hd__dfxtp_1
X_15084_ _07128_ _07207_ _07206_ vssd1 vssd1 vccd1 vccd1 _07772_ sky130_fd_sc_hd__a21oi_1
XFILLER_181_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12296_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] _05052_
+ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__a21o_1
XFILLER_10_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14035_ _06773_ vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__clkbuf_1
X_11247_ gpout0.hpos\[2\] gpout0.hpos\[1\] vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__nand2_1
XFILLER_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19892_ clknet_leaf_14_i_clk _00823_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18843_ rbzero.debug_overlay.vplaneY\[-6\] _02634_ vssd1 vssd1 vccd1 vccd1 _02684_
+ sky130_fd_sc_hd__and2_1
X_11178_ rbzero.tex_r1\[2\] _03926_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__or2_1
XFILLER_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10129_ _03122_ vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__clkbuf_1
X_18774_ rbzero.pov.ready_buffer\[37\] _02644_ _02646_ _02559_ vssd1 vssd1 vccd1 vccd1
+ _01030_ sky130_fd_sc_hd__a211o_1
X_15986_ _07269_ _08333_ _08332_ _08330_ vssd1 vssd1 vccd1 vccd1 _08600_ sky130_fd_sc_hd__o31a_1
XFILLER_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17725_ _01980_ _01991_ _01995_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__o21a_1
X_14937_ _06978_ _07006_ _07157_ _07178_ vssd1 vssd1 vccd1 vccd1 _07625_ sky130_fd_sc_hd__or4_1
XFILLER_94_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18929__114 clknet_1_1__leaf__02724_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__inv_2
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17656_ _01932_ vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14868_ _06977_ _07147_ _07554_ _07555_ vssd1 vssd1 vccd1 vccd1 _07556_ sky130_fd_sc_hd__or4_1
XFILLER_91_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16607_ _08643_ _07960_ _09215_ vssd1 vssd1 vccd1 vccd1 _09216_ sky130_fd_sc_hd__or3b_1
X_13819_ _05616_ _06056_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__nor2_1
XFILLER_90_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17587_ _01786_ _01757_ _01872_ vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__a21oi_1
XFILLER_189_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14799_ _07481_ _07486_ vssd1 vssd1 vccd1 vccd1 _07487_ sky130_fd_sc_hd__or2b_1
XFILLER_50_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19326_ rbzero.traced_texa\[0\] rbzero.texV\[0\] vssd1 vssd1 vccd1 vccd1 _02812_
+ sky130_fd_sc_hd__nand2_1
X_16538_ _09146_ _09147_ vssd1 vssd1 vccd1 vccd1 _09148_ sky130_fd_sc_hd__and2b_1
X_19257_ gpout5.clk_div\[0\] net61 vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__nor2_1
X_16469_ _09076_ _09079_ _08485_ vssd1 vssd1 vccd1 vccd1 _09080_ sky130_fd_sc_hd__o21ai_1
X_18208_ rbzero.color_sky\[2\] rbzero.spi_registers.new_sky\[2\] _02320_ vssd1 vssd1
+ vccd1 vccd1 _02326_ sky130_fd_sc_hd__mux2_1
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18139_ _02281_ _03902_ _02258_ vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__or3b_1
XFILLER_172_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18975__156 clknet_1_1__leaf__02728_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__inv_2
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20101_ clknet_leaf_88_i_clk _01032_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
X_09912_ _03008_ vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20032_ clknet_leaf_86_i_clk _00963_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_09843_ _02970_ vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__clkbuf_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09774_ _02934_ vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_60_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19047__220 clknet_1_1__leaf__02736_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__inv_2
XFILLER_170_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_75_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_41_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10480_ _03306_ vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19093__262 clknet_1_0__leaf__02740_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__inv_2
X_12150_ _04876_ _04874_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__nand2_1
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11101_ _03860_ _03868_ _03886_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_13_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12081_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] vssd1
+ vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__nand2_1
X_11032_ _02902_ _03797_ _03799_ _03817_ _02903_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__o221a_1
XFILLER_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15840_ rbzero.map_rom.i_col\[4\] _07825_ vssd1 vssd1 vccd1 vccd1 _08470_ sky130_fd_sc_hd__nor2_1
XFILLER_77_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _08443_ _08439_ _08444_ vssd1 vssd1 vccd1 vccd1 _08445_ sky130_fd_sc_hd__and3b_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ _05707_ _05734_ _05739_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__a21o_1
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17510_ _01797_ _01798_ _01799_ _01800_ vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__a211o_1
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14722_ _06865_ _07039_ vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__or2_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18490_ rbzero.pov.spi_buffer\[15\] rbzero.pov.spi_buffer\[16\] _02455_ vssd1 vssd1
+ vccd1 vccd1 _02462_ sky130_fd_sc_hd__mux2_1
X_11934_ net25 vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__inv_2
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ rbzero.debug_overlay.vplaneY\[-3\] rbzero.wall_tracer.rayAddendY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__nand2_1
XFILLER_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14653_ _07308_ _07315_ vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__xnor2_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ net51 _04625_ _04626_ net53 vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__a22o_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _06319_ _06318_ _06312_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__a21o_1
X_10816_ _03570_ _03601_ rbzero.row_render.vinf vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__a21oi_1
X_17372_ _01678_ vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14584_ _07268_ _07271_ vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__xnor2_1
X_11796_ net47 _04569_ _04570_ _04572_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__a22o_1
XFILLER_14_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16323_ _08932_ _08934_ vssd1 vssd1 vccd1 vccd1 _08935_ sky130_fd_sc_hd__nor2_1
X_13535_ _06289_ _06290_ vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__nand2_1
XFILLER_186_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10747_ gpout0.vpos\[9\] _03469_ net1 vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__or3b_1
XFILLER_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16254_ _07735_ _07333_ _08865_ vssd1 vssd1 vccd1 vccd1 _08866_ sky130_fd_sc_hd__or3_1
XFILLER_158_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13466_ _06219_ _06221_ vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__nand2_1
X_10678_ gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__inv_2
XFILLER_174_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15205_ _07673_ _07173_ vssd1 vssd1 vccd1 vccd1 _07892_ sky130_fd_sc_hd__nand2_1
X_12417_ _05170_ _05172_ _05173_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__mux2_1
X_16185_ _07877_ _08018_ vssd1 vssd1 vccd1 vccd1 _08798_ sky130_fd_sc_hd__nor2_1
X_13397_ _06147_ _06153_ _06145_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__o21ba_1
XFILLER_142_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15136_ _07822_ _07823_ vssd1 vssd1 vccd1 vccd1 _07824_ sky130_fd_sc_hd__nand2_1
XFILLER_182_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12348_ _03487_ _05102_ _05103_ _05104_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__a22o_2
XFILLER_99_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19944_ net173 _00875_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[24\] sky130_fd_sc_hd__dfxtp_1
X_15067_ _07178_ _07176_ _07754_ vssd1 vssd1 vccd1 vccd1 _07755_ sky130_fd_sc_hd__or3_1
X_12279_ rbzero.debug_overlay.facingX\[-5\] rbzero.wall_tracer.rayAddendX\[3\] vssd1
+ vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__or2_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14018_ rbzero.wall_tracer.stepDistY\[4\] _06759_ _06718_ vssd1 vssd1 vccd1 vccd1
+ _06760_ sky130_fd_sc_hd__mux2_1
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19875_ clknet_leaf_22_i_clk _00806_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18826_ rbzero.pov.ready_buffer\[16\] _02666_ _02674_ _02675_ vssd1 vssd1 vccd1 vccd1
+ _01053_ sky130_fd_sc_hd__a211o_1
XFILLER_95_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18757_ _02633_ vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__buf_2
XFILLER_49_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15969_ _04946_ _08431_ vssd1 vssd1 vccd1 vccd1 _08584_ sky130_fd_sc_hd__nand2_1
X_17708_ _04100_ _01959_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__nor2_1
XFILLER_36_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18688_ _02578_ _02580_ _02266_ vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__o21a_1
XFILLER_64_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17639_ rbzero.debug_overlay.vplaneX\[-5\] rbzero.wall_tracer.rayAddendX\[-5\] vssd1
+ vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__nor2_1
XFILLER_36_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19309_ _02794_ _02795_ _02797_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__or3_1
XFILLER_149_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20015_ clknet_leaf_92_i_clk _00946_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_09826_ _02961_ vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_115_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09757_ _02925_ vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11650_ _03607_ _04426_ _04430_ _03704_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__a211o_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10601_ _03346_ _03375_ _03359_ _03391_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__nor4_1
XFILLER_70_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11581_ rbzero.tex_b0\[25\] rbzero.tex_b0\[24\] _04189_ vssd1 vssd1 vccd1 vccd1 _04363_
+ sky130_fd_sc_hd__mux2_1
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10532_ _03333_ vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__clkbuf_1
X_13320_ _06000_ _06067_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__xor2_1
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10463_ _03297_ vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__clkbuf_1
X_13251_ _05474_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__clkbuf_4
XFILLER_108_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18958__140 clknet_1_0__leaf__02727_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__inv_2
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12202_ rbzero.wall_tracer.trackDistY\[-1\] vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__inv_2
X_13182_ _05910_ _05938_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__or2b_1
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10394_ _03261_ vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12133_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__or2_1
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17990_ rbzero.pov.spi_buffer\[48\] rbzero.pov.ready_buffer\[48\] _02186_ vssd1 vssd1
+ vccd1 vccd1 _02196_ sky130_fd_sc_hd__mux2_1
XFILLER_97_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16941_ _09016_ _09546_ vssd1 vssd1 vccd1 vccd1 _09547_ sky130_fd_sc_hd__or2_1
X_12064_ net72 rbzero.wall_tracer.state\[4\] _02907_ vssd1 vssd1 vccd1 vccd1 _04833_
+ sky130_fd_sc_hd__and3_2
XFILLER_78_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11015_ _03775_ _03800_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__nor2_1
X_19660_ clknet_leaf_15_i_clk _00591_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16872_ _09384_ _09376_ vssd1 vssd1 vccd1 vccd1 _09479_ sky130_fd_sc_hd__or2b_1
XFILLER_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18611_ _04532_ rbzero.pov.mosi_buffer\[0\] _03337_ vssd1 vssd1 vccd1 vccd1 _02525_
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15823_ rbzero.traced_texa\[3\] _08461_ _08462_ rbzero.wall_tracer.visualWallDist\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__a22o_1
XFILLER_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19591_ clknet_leaf_40_i_clk _00522_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18542_ _02489_ vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__clkbuf_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ rbzero.wall_tracer.texu\[5\] _06853_ _08435_ _08436_ _03485_ vssd1 vssd1
+ vccd1 vccd1 _00480_ sky130_fd_sc_hd__o221a_1
X_12966_ _05664_ _05681_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__or2_1
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14705_ _07376_ _07392_ vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__xnor2_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18473_ rbzero.pov.spi_buffer\[7\] rbzero.pov.spi_buffer\[8\] _02444_ vssd1 vssd1
+ vccd1 vccd1 _02453_ sky130_fd_sc_hd__mux2_1
X_11917_ _03906_ _04499_ _03909_ _04500_ _04691_ _04672_ vssd1 vssd1 vccd1 vccd1 _04692_
+ sky130_fd_sc_hd__mux4_1
X_15685_ _07494_ _08252_ _07766_ _06997_ vssd1 vssd1 vccd1 vccd1 _08368_ sky130_fd_sc_hd__o22ai_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _05505_ _05502_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__nor2_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17424_ _03340_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__clkbuf_4
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _07312_ _07320_ _07322_ vssd1 vssd1 vccd1 vccd1 _07324_ sky130_fd_sc_hd__nand3_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ net11 vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__inv_2
XFILLER_21_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17355_ rbzero.spi_registers.new_mapd\[6\] rbzero.spi_registers.spi_buffer\[6\] _01663_
+ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__mux2_1
X_14567_ _07253_ _07254_ vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__nand2_1
XFILLER_147_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11779_ _04552_ net62 vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__or2_1
XFILLER_119_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16306_ _08910_ _08916_ vssd1 vssd1 vccd1 vccd1 _08918_ sky130_fd_sc_hd__or2_1
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13518_ _06232_ _06234_ _06252_ _06274_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__a31o_1
X_17286_ _01534_ _01613_ _01614_ _01526_ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__a31o_1
XFILLER_201_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14498_ _07154_ _07185_ _07179_ vssd1 vssd1 vccd1 vccd1 _07186_ sky130_fd_sc_hd__or3_1
XFILLER_158_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16237_ _07972_ _08191_ vssd1 vssd1 vccd1 vccd1 _08849_ sky130_fd_sc_hd__nor2_1
X_13449_ _06116_ _06138_ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__nor2_1
XFILLER_162_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16168_ _08779_ _08780_ vssd1 vssd1 vccd1 vccd1 _08781_ sky130_fd_sc_hd__nor2_1
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15119_ _07805_ _07806_ vssd1 vssd1 vccd1 vccd1 _07807_ sky130_fd_sc_hd__xnor2_4
XFILLER_138_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16099_ _08711_ _08712_ vssd1 vssd1 vccd1 vccd1 _08713_ sky130_fd_sc_hd__nand2_2
XFILLER_86_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19927_ net156 _00858_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19230__386 clknet_1_0__leaf__02753_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__inv_2
XFILLER_96_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19858_ clknet_leaf_23_i_clk _00789_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18809_ rbzero.pov.ready_buffer\[31\] _02644_ _02665_ _02651_ vssd1 vssd1 vccd1 vccd1
+ _01046_ sky130_fd_sc_hd__a211o_1
X_19789_ clknet_leaf_87_i_clk _00720_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19159__321 clknet_1_0__leaf__02747_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__inv_2
XFILLER_165_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20495_ clknet_leaf_43_i_clk _01426_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09809_ _02952_ vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12820_ _05491_ _05576_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__nand2_1
XFILLER_27_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _05467_ _05483_ _05473_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__a21oi_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _03783_ _02899_ _04236_ _04481_ _03527_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__a311o_1
X_15470_ _08129_ _08026_ _08153_ vssd1 vssd1 vccd1 vccd1 _08155_ sky130_fd_sc_hd__and3_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _05436_ _05438_ _05333_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__a21o_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14421_ _04949_ _07102_ _07107_ _07108_ vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__a22o_1
X_11633_ _03674_ _04413_ _03704_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__a21o_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17140_ _09133_ _07961_ vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__nor2_1
XFILLER_168_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14352_ _06978_ _07037_ vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__or2_1
XFILLER_196_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11564_ _03656_ _04343_ _04344_ _04345_ _03606_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__o221a_1
XFILLER_129_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13303_ _05480_ _06056_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__nand2_2
X_17071_ _09231_ _09256_ _09229_ _09142_ vssd1 vssd1 vccd1 vccd1 _09676_ sky130_fd_sc_hd__o22a_1
X_10515_ rbzero.tex_b0\[12\] rbzero.tex_b0\[11\] _03324_ vssd1 vssd1 vccd1 vccd1 _03325_
+ sky130_fd_sc_hd__mux2_1
X_11495_ rbzero.tex_g1\[55\] rbzero.tex_g1\[54\] _03617_ vssd1 vssd1 vccd1 vccd1 _04278_
+ sky130_fd_sc_hd__mux2_1
X_14283_ _06940_ _06968_ _06969_ _06970_ vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__o22ai_1
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16022_ _08604_ _08635_ vssd1 vssd1 vccd1 vccd1 _08636_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10446_ _03288_ vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__clkbuf_1
X_13234_ _05906_ _05949_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10377_ _03252_ vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13165_ _05870_ _05920_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__nand2_1
XFILLER_123_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12116_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[9\] vssd1
+ vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__and2_1
XFILLER_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17973_ _02187_ vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__clkbuf_1
X_13096_ _05761_ _05763_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__nor2_1
XFILLER_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16924_ _09527_ _09462_ _09528_ vssd1 vssd1 vccd1 vccd1 _09530_ sky130_fd_sc_hd__and3_1
X_12047_ net50 net51 net53 _04532_ _04779_ net34 vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__mux4_1
X_19712_ clknet_leaf_2_i_clk _00643_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16855_ _09460_ _09461_ vssd1 vssd1 vccd1 vccd1 _09462_ sky130_fd_sc_hd__or2b_1
X_19643_ clknet_leaf_51_i_clk _00574_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15806_ _08452_ vssd1 vssd1 vccd1 vccd1 _08458_ sky130_fd_sc_hd__buf_4
XFILLER_92_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19574_ clknet_leaf_41_i_clk _00505_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_16786_ _09267_ _09288_ _09286_ vssd1 vssd1 vccd1 vccd1 _09394_ sky130_fd_sc_hd__a21oi_2
XFILLER_168_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13998_ _05315_ _06714_ _06741_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__o21ai_1
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18525_ _02480_ vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__clkbuf_1
X_15737_ _08355_ _08419_ vssd1 vssd1 vccd1 vccd1 _08420_ sky130_fd_sc_hd__xnor2_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12949_ _05465_ _05697_ _05479_ _05538_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__a22o_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18456_ _02443_ vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__clkbuf_4
XFILLER_61_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15668_ _08335_ _08350_ vssd1 vssd1 vccd1 vccd1 _08351_ sky130_fd_sc_hd__xnor2_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17407_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.wall_tracer.rayAddendY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__nor2_1
XFILLER_92_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14619_ _07301_ _07305_ _07306_ vssd1 vssd1 vccd1 vccd1 _07307_ sky130_fd_sc_hd__a21bo_1
XFILLER_60_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15599_ _08281_ _08282_ vssd1 vssd1 vccd1 vccd1 _08283_ sky130_fd_sc_hd__xor2_1
XFILLER_21_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17338_ rbzero.spi_registers.spi_cmd\[0\] _01658_ rbzero.spi_registers.spi_cmd\[3\]
+ rbzero.spi_registers.spi_cmd\[2\] vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__or4b_2
XFILLER_186_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17269_ _01595_ _01596_ _01597_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__a21o_1
XFILLER_140_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20280_ net340 _01211_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10300_ _03212_ vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11280_ _03463_ _04040_ _04052_ _04062_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__or4b_2
XFILLER_153_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20478_ clknet_leaf_66_i_clk _01409_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10231_ rbzero.tex_g0\[19\] rbzero.tex_g0\[18\] _03166_ vssd1 vssd1 vccd1 vccd1 _03176_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10162_ _03139_ vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19213__370 clknet_1_0__leaf__02752_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__inv_2
XFILLER_120_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10093_ _03103_ vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__clkbuf_1
X_14970_ _07656_ _07657_ vssd1 vssd1 vccd1 vccd1 _07658_ sky130_fd_sc_hd__nor2_1
XFILLER_0_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13921_ _05333_ _06673_ _05369_ vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__a21oi_1
XFILLER_101_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16640_ _07012_ _08130_ _07173_ _08766_ vssd1 vssd1 vccd1 vccd1 _09249_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_142_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13852_ _06435_ _06608_ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__xor2_2
XFILLER_47_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12803_ _05558_ _05559_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__nand2_1
XFILLER_76_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16571_ _09130_ _09180_ vssd1 vssd1 vccd1 vccd1 _09181_ sky130_fd_sc_hd__xnor2_1
X_13783_ _06515_ _06528_ vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__xor2_1
X_10995_ gpout0.hpos\[5\] vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__inv_2
XFILLER_71_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18310_ _02389_ vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15522_ _07235_ _07786_ vssd1 vssd1 vccd1 vccd1 _08206_ sky130_fd_sc_hd__nor2_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12734_ _05465_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__buf_2
X_19290_ rbzero.traced_texa\[-6\] rbzero.texV\[-6\] vssd1 vssd1 vccd1 vccd1 _02782_
+ sky130_fd_sc_hd__xnor2_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ rbzero.spi_registers.got_new_vshift _02262_ vssd1 vssd1 vccd1 vccd1 _02349_
+ sky130_fd_sc_hd__and2_1
XFILLER_188_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15453_ _07213_ _07897_ vssd1 vssd1 vccd1 vccd1 _08138_ sky130_fd_sc_hd__nor2_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12665_ _05421_ _05396_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__or2_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _07091_ vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__clkbuf_4
XFILLER_169_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11616_ rbzero.row_render.texu\[0\] _03729_ _03730_ _03996_ vssd1 vssd1 vccd1 vccd1
+ _04397_ sky130_fd_sc_hd__a31o_1
X_18172_ rbzero.map_overlay.i_mapdy\[4\] _02291_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__or2_1
X_15384_ rbzero.wall_tracer.visualWallDist\[8\] _07256_ vssd1 vssd1 vccd1 vccd1 _08069_
+ sky130_fd_sc_hd__nand2_1
X_12596_ _05310_ _05332_ _05335_ _05352_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__a31o_1
XFILLER_129_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17123_ _08899_ _08333_ vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__nor2_1
XFILLER_7_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14335_ _07021_ _07022_ _06914_ vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__mux2_1
X_11547_ rbzero.tex_b0\[54\] _04247_ _03652_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__a21o_1
XFILLER_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17054_ _09559_ _09537_ vssd1 vssd1 vccd1 vccd1 _09659_ sky130_fd_sc_hd__or2b_1
X_14266_ _04838_ rbzero.wall_tracer.stepDistX\[-6\] _06950_ _06953_ vssd1 vssd1 vccd1
+ vccd1 _06954_ sky130_fd_sc_hd__o22ai_4
X_11478_ rbzero.tex_g1\[11\] rbzero.tex_g1\[10\] _03618_ vssd1 vssd1 vccd1 vccd1 _04261_
+ sky130_fd_sc_hd__mux2_1
XFILLER_171_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16005_ _07097_ _07084_ _07332_ _07786_ vssd1 vssd1 vccd1 vccd1 _08619_ sky130_fd_sc_hd__or4_1
Xclkbuf_0__02743_ _02743_ vssd1 vssd1 vccd1 vccd1 clknet_0__02743_ sky130_fd_sc_hd__clkbuf_16
X_13217_ _05972_ _05973_ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__nor2_1
X_10429_ _03279_ vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14197_ _05137_ _05086_ _05143_ _06884_ vssd1 vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__and4b_1
XFILLER_140_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _05901_ _05904_ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__nor2_1
XFILLER_98_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _05801_ _05835_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__xor2_2
X_17956_ _02178_ vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16907_ _09318_ _09513_ vssd1 vssd1 vccd1 vccd1 _09514_ sky130_fd_sc_hd__xnor2_1
X_17887_ rbzero.pov.spi_done _02907_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__nand2_1
XFILLER_65_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19626_ clknet_leaf_45_i_clk _00557_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16838_ _09358_ _09360_ _09357_ vssd1 vssd1 vccd1 vccd1 _09445_ sky130_fd_sc_hd__a21bo_1
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16769_ _08247_ _07530_ _08681_ vssd1 vssd1 vccd1 vccd1 _09377_ sky130_fd_sc_hd__or3_1
XFILLER_19_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19557_ clknet_leaf_11_i_clk _00488_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18508_ _02471_ vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19488_ clknet_leaf_52_i_clk _00434_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19041__215 clknet_1_0__leaf__02735_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__inv_2
XFILLER_22_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20401_ net461 _01332_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20332_ net392 _01263_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20263_ net323 _01194_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20194_ net254 _01125_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02732_ clknet_0__02732_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02732_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_99_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _03565_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__inv_2
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ _05202_ _05203_ _05204_ _05206_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__a211oi_2
XFILLER_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11401_ _03704_ _04175_ _04180_ _04184_ _03684_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__o221a_1
XFILLER_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12381_ _05072_ _05137_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__or2_1
XFILLER_153_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14120_ _06824_ vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_193_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11332_ rbzero.debug_overlay.facingX\[-6\] _04084_ _03901_ gpout0.vpos\[5\] vssd1
+ vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__a211o_1
XFILLER_197_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14051_ _06785_ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__clkbuf_4
X_11263_ _04037_ _04047_ _03513_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__o21ba_1
XFILLER_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13002_ _05732_ _05757_ _05758_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10214_ _03167_ vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11194_ rbzero.tex_r1\[29\] _03660_ _03768_ _03702_ vssd1 vssd1 vccd1 vccd1 _03979_
+ sky130_fd_sc_hd__a31o_1
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10145_ _03130_ vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__clkbuf_1
X_17810_ _02072_ _02073_ _02068_ _02069_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__a211o_1
X_18790_ rbzero.debug_overlay.facingY\[-8\] _02638_ vssd1 vssd1 vccd1 vccd1 _02655_
+ sky130_fd_sc_hd__or2_1
XFILLER_43_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17741_ rbzero.wall_tracer.rayAddendX\[2\] rbzero.wall_tracer.rayAddendX\[1\] _01985_
+ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__o21ai_1
X_10076_ _03094_ vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__clkbuf_1
X_14953_ _07575_ _07612_ _07613_ _07640_ vssd1 vssd1 vccd1 vccd1 _07641_ sky130_fd_sc_hd__and4_1
XFILLER_48_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13904_ rbzero.wall_tracer.stepDistY\[-9\] _06658_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _06659_ sky130_fd_sc_hd__mux2_1
X_17672_ _01942_ _01943_ _01945_ _01946_ _03497_ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__o311a_1
XFILLER_78_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14884_ _07480_ _07524_ vssd1 vssd1 vccd1 vccd1 _07572_ sky130_fd_sc_hd__xor2_1
X_16623_ _08252_ _09231_ vssd1 vssd1 vccd1 vccd1 _09232_ sky130_fd_sc_hd__nor2_1
X_19411_ _08452_ _01705_ _02872_ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__and3_1
XFILLER_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13835_ _06577_ _06590_ _06591_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__a21oi_2
XFILLER_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16554_ _09154_ _09163_ vssd1 vssd1 vccd1 vccd1 _09164_ sky130_fd_sc_hd__xor2_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19342_ _02825_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__inv_2
X_13766_ _06518_ _06522_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10978_ net41 vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__inv_2
XFILLER_43_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15505_ _08114_ _08094_ vssd1 vssd1 vccd1 vccd1 _08189_ sky130_fd_sc_hd__or2b_1
XFILLER_188_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12717_ _05392_ _05467_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__xor2_4
X_19273_ rbzero.traced_texa\[-9\] rbzero.texV\[-9\] vssd1 vssd1 vccd1 vccd1 _02768_
+ sky130_fd_sc_hd__nor2_1
X_16485_ _09002_ _09093_ _09094_ vssd1 vssd1 vccd1 vccd1 _09095_ sky130_fd_sc_hd__a21oi_2
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13697_ _05805_ _05992_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__nor2_1
XFILLER_70_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18224_ _02337_ vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__clkbuf_1
X_15436_ _06997_ _07138_ vssd1 vssd1 vccd1 vccd1 _08121_ sky130_fd_sc_hd__nor2_1
X_12648_ _05256_ _05228_ _05313_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__mux2_1
XFILLER_54_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18155_ rbzero.map_overlay.i_mapdx\[2\] _02292_ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__or2_1
XFILLER_200_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15367_ rbzero.debug_overlay.playerY\[-4\] rbzero.debug_overlay.playerX\[-4\] _06851_
+ vssd1 vssd1 vccd1 vccd1 _08053_ sky130_fd_sc_hd__mux2_1
XFILLER_102_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12579_ _05305_ _05302_ _05306_ _05189_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__or4b_1
XFILLER_157_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17106_ rbzero.wall_tracer.trackDistX\[9\] rbzero.wall_tracer.stepDistX\[9\] vssd1
+ vssd1 vccd1 vccd1 _09711_ sky130_fd_sc_hd__or2_1
X_14318_ _07005_ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__buf_2
XFILLER_50_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18086_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[2\] _02245_
+ vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__mux2_1
XFILLER_116_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15298_ _07084_ vssd1 vssd1 vccd1 vccd1 _07984_ sky130_fd_sc_hd__clkbuf_4
XFILLER_7_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17037_ _09014_ _09016_ _08803_ vssd1 vssd1 vccd1 vccd1 _09642_ sky130_fd_sc_hd__a21oi_1
X_14249_ _06852_ _06695_ _06936_ _06859_ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__o211a_1
XFILLER_125_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__02726_ _02726_ vssd1 vssd1 vccd1 vccd1 clknet_0__02726_ sky130_fd_sc_hd__clkbuf_16
XFILLER_98_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _02942_ vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__clkbuf_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ _02169_ vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19609_ clknet_leaf_55_i_clk _00540_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20315_ net375 _01246_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20246_ net306 _01177_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18952__135 clknet_1_1__leaf__02726_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__inv_2
XFILLER_131_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20177_ net237 _01108_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09988_ rbzero.tex_r0\[6\] rbzero.tex_r0\[5\] _03039_ vssd1 vssd1 vccd1 vccd1 _03048_
+ sky130_fd_sc_hd__mux2_1
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ net28 net27 vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__nor2_1
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ _03603_ _03683_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__nor2_4
Xtop_ew_algofoogle_108 vssd1 vssd1 vccd1 vccd1 ones[1] top_ew_algofoogle_108/LO sky130_fd_sc_hd__conb_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtop_ew_algofoogle_119 vssd1 vssd1 vccd1 vccd1 ones[12] top_ew_algofoogle_119/LO sky130_fd_sc_hd__conb_1
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11881_ net10 _04656_ _04645_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__o21ai_1
XFILLER_45_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13620_ _06359_ _06375_ _06376_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__a21boi_1
XFILLER_72_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10832_ _03617_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__buf_4
XFILLER_72_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13551_ _06255_ _06267_ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10763_ rbzero.texV\[3\] _03547_ _03548_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a21boi_2
XFILLER_186_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12502_ _05225_ _05258_ _05247_ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__or3_1
X_16270_ _08847_ _08881_ vssd1 vssd1 vccd1 vccd1 _08882_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13482_ _06143_ _06238_ vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__xor2_1
XFILLER_157_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10694_ _03480_ _03481_ _03482_ _03485_ _00000_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__a41o_1
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15221_ _07746_ _07763_ _07907_ vssd1 vssd1 vccd1 vccd1 _07908_ sky130_fd_sc_hd__a21oi_2
XFILLER_157_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12433_ _05138_ _05140_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__nand2_1
XFILLER_200_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15152_ rbzero.wall_tracer.visualWallDist\[6\] _07256_ vssd1 vssd1 vccd1 vccd1 _07839_
+ sky130_fd_sc_hd__nand2_1
X_12364_ _05040_ _05041_ _05042_ vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__o21a_1
XFILLER_138_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14103_ rbzero.wall_tracer.stepDistX\[-11\] _06631_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _06816_ sky130_fd_sc_hd__mux2_1
XFILLER_181_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11315_ rbzero.debug_overlay.vplaneX\[-5\] vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__clkbuf_4
XFILLER_5_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19960_ net189 _00891_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15083_ _07741_ _07770_ vssd1 vssd1 vccd1 vccd1 _07771_ sky130_fd_sc_hd__xnor2_1
X_12295_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] vssd1
+ vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__or2_1
XFILLER_99_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14034_ rbzero.wall_tracer.stepDistY\[7\] _06772_ _06718_ vssd1 vssd1 vccd1 vccd1
+ _06773_ sky130_fd_sc_hd__mux2_1
XFILLER_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11246_ _03896_ _04004_ _04030_ _03897_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__o2bb2a_1
X_19891_ clknet_leaf_21_i_clk _00822_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_leak
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19070__241 clknet_1_0__leaf__02738_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__inv_2
X_18842_ rbzero.pov.ready_buffer\[2\] _02635_ _02683_ _02672_ vssd1 vssd1 vccd1 vccd1
+ _01061_ sky130_fd_sc_hd__o211a_1
XFILLER_164_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11177_ rbzero.tex_r1\[4\] _03661_ _03936_ _03961_ vssd1 vssd1 vccd1 vccd1 _03962_
+ sky130_fd_sc_hd__a31o_1
XFILLER_68_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10128_ rbzero.tex_g1\[3\] rbzero.tex_g1\[4\] _03117_ vssd1 vssd1 vccd1 vccd1 _03122_
+ sky130_fd_sc_hd__mux2_1
X_15985_ _08354_ _08323_ vssd1 vssd1 vccd1 vccd1 _08599_ sky130_fd_sc_hd__or2b_1
X_18773_ rbzero.debug_overlay.facingX\[-5\] _02645_ vssd1 vssd1 vccd1 vccd1 _02646_
+ sky130_fd_sc_hd__and2_1
XFILLER_95_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14936_ _06979_ _07185_ _07199_ _07006_ vssd1 vssd1 vccd1 vccd1 _07624_ sky130_fd_sc_hd__o22a_1
X_10059_ rbzero.tex_g1\[36\] rbzero.tex_g1\[37\] _03084_ vssd1 vssd1 vccd1 vccd1 _03086_
+ sky130_fd_sc_hd__mux2_1
X_17724_ _01977_ _01994_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17655_ rbzero.wall_tracer.rayAddendX\[-5\] _01931_ _03509_ vssd1 vssd1 vccd1 vccd1
+ _01932_ sky130_fd_sc_hd__mux2_1
X_14867_ _06938_ _07156_ _07177_ _06954_ vssd1 vssd1 vccd1 vccd1 _07555_ sky130_fd_sc_hd__o22a_1
XFILLER_24_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16606_ _07123_ _08070_ vssd1 vssd1 vccd1 vccd1 _09215_ sky130_fd_sc_hd__nor2_1
XFILLER_51_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13818_ _06227_ _06570_ _06574_ _06211_ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__a22o_1
XFILLER_91_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17586_ _01757_ rbzero.debug_overlay.vplaneY\[-1\] _01785_ vssd1 vssd1 vccd1 vccd1
+ _01872_ sky130_fd_sc_hd__a21oi_1
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14798_ _06933_ _07006_ _07485_ _07484_ vssd1 vssd1 vccd1 vccd1 _07486_ sky130_fd_sc_hd__o31ai_1
XFILLER_90_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16537_ _09144_ _09145_ vssd1 vssd1 vccd1 vccd1 _09147_ sky130_fd_sc_hd__nand2_1
X_19325_ rbzero.traced_texa\[0\] rbzero.texV\[0\] vssd1 vssd1 vccd1 vccd1 _02811_
+ sky130_fd_sc_hd__or2_1
XFILLER_188_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13749_ _06478_ _06505_ vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__xor2_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16468_ _09077_ _08957_ _09078_ vssd1 vssd1 vccd1 vccd1 _09079_ sky130_fd_sc_hd__a21oi_2
XFILLER_32_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15419_ _07979_ _08102_ _08103_ vssd1 vssd1 vccd1 vccd1 _08104_ sky130_fd_sc_hd__a21bo_1
X_18207_ _02325_ vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__clkbuf_1
X_19187_ clknet_1_0__leaf__02743_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__buf_1
X_16399_ _09007_ _08899_ _08896_ _09009_ vssd1 vssd1 vccd1 vccd1 _09010_ sky130_fd_sc_hd__o22ai_1
XFILLER_157_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18138_ _04503_ _02280_ vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__nand2_1
XFILLER_191_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19153__316 clknet_1_0__leaf__02746_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__inv_2
X_18069_ _02238_ vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__clkbuf_1
XFILLER_105_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20100_ clknet_leaf_88_i_clk _01031_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_176_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09911_ rbzero.tex_r0\[43\] rbzero.tex_r0\[42\] _03006_ vssd1 vssd1 vccd1 vccd1 _03008_
+ sky130_fd_sc_hd__mux2_1
XFILLER_160_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20031_ clknet_leaf_85_i_clk _00962_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09842_ rbzero.tex_r1\[9\] rbzero.tex_r1\[10\] _02965_ vssd1 vssd1 vccd1 vccd1 _02970_
+ sky130_fd_sc_hd__mux2_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ rbzero.tex_r1\[42\] rbzero.tex_r1\[43\] _02932_ vssd1 vssd1 vccd1 vccd1 _02934_
+ sky130_fd_sc_hd__mux2_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_9_i_clk clknet_opt_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18388__32 clknet_1_0__leaf__02434_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__inv_2
XFILLER_15_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11100_ _03870_ _03878_ _03885_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__or3_1
XFILLER_123_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12080_ _04842_ vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11031_ _03466_ _03801_ _03798_ _02900_ _03816_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__o221a_1
X_20229_ net289 _01160_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_49_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15770_ _02901_ _03838_ _04034_ _03459_ vssd1 vssd1 vccd1 vccd1 _08444_ sky130_fd_sc_hd__a31o_1
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _05735_ _05736_ _05738_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__a21bo_1
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14721_ _07375_ _07408_ vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__xor2_1
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11933_ net22 _04670_ _04680_ _04707_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__and4_1
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17440_ _04109_ rbzero.wall_tracer.rayAddendY\[-2\] vssd1 vssd1 vccd1 vccd1 _01736_
+ sky130_fd_sc_hd__and2_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _07318_ _07326_ vssd1 vssd1 vccd1 vccd1 _07340_ sky130_fd_sc_hd__xnor2_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ gpout1.clk_div\[1\] _04627_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__or2b_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _06319_ _06312_ _06318_ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__nand3_1
XFILLER_72_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _03576_ _03582_ _03599_ _03600_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__o31a_1
X_17371_ rbzero.spi_registers.new_mapd\[14\] rbzero.spi_registers.spi_buffer\[14\]
+ _01662_ vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__mux2_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ _07269_ _07270_ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__nor2_1
X_11795_ _04532_ _04571_ net48 vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__a21o_1
X_16322_ _08797_ _08811_ _08933_ vssd1 vssd1 vccd1 vccd1 _08934_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13534_ _06289_ _06290_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__xnor2_1
X_10746_ _03517_ _03518_ _03531_ gpout0.vpos\[8\] vssd1 vssd1 vccd1 vccd1 _03532_
+ sky130_fd_sc_hd__o31a_1
XFILLER_199_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16253_ _07123_ _07787_ vssd1 vssd1 vccd1 vccd1 _08865_ sky130_fd_sc_hd__or2_1
XFILLER_158_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13465_ _06219_ _06221_ vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__or2_1
XFILLER_159_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10677_ _03461_ _03465_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__nor2_1
X_15204_ _07887_ _07890_ vssd1 vssd1 vccd1 vccd1 _07891_ sky130_fd_sc_hd__xor2_2
XFILLER_51_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12416_ _05077_ _05150_ _05166_ _05152_ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__a31o_1
XFILLER_199_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16184_ _08787_ _08796_ vssd1 vssd1 vccd1 vccd1 _08797_ sky130_fd_sc_hd__xor2_2
XFILLER_166_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13396_ _06001_ _05988_ _06148_ _06152_ vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__o31a_1
XFILLER_182_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15135_ _07812_ _07821_ vssd1 vssd1 vccd1 vccd1 _07823_ sky130_fd_sc_hd__nand2_1
X_12347_ rbzero.wall_tracer.visualWallDist\[-6\] _03479_ _05072_ vssd1 vssd1 vccd1
+ vccd1 _05104_ sky130_fd_sc_hd__o21a_1
XFILLER_181_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19943_ net172 _00874_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[23\] sky130_fd_sc_hd__dfxtp_1
X_15066_ _04840_ rbzero.wall_tracer.stepDistX\[5\] _07752_ _07753_ vssd1 vssd1 vccd1
+ vccd1 _07754_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12278_ rbzero.debug_overlay.facingX\[-5\] rbzero.wall_tracer.rayAddendX\[3\] vssd1
+ vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__nand2_1
XFILLER_49_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14017_ _06758_ vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__buf_2
XFILLER_68_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11229_ gpout0.vpos\[4\] _03524_ _03523_ gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1
+ _04014_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19874_ clknet_leaf_22_i_clk _00805_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18825_ _03338_ vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__buf_4
XFILLER_56_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18756_ _02288_ _02632_ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__nand2_1
X_15968_ rbzero.wall_tracer.trackDistX\[-2\] _08553_ _08577_ _08583_ vssd1 vssd1 vccd1
+ vccd1 _00547_ sky130_fd_sc_hd__o22a_1
XFILLER_76_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17707_ _01977_ _01978_ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__nand2_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14919_ _07605_ _07606_ vssd1 vssd1 vccd1 vccd1 _07607_ sky130_fd_sc_hd__and2_1
XFILLER_64_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18687_ rbzero.pov.ready_buffer\[73\] _02540_ _02543_ _02579_ vssd1 vssd1 vccd1 vccd1
+ _02580_ sky130_fd_sc_hd__o211a_1
X_15899_ _08512_ _08520_ _08521_ _08522_ vssd1 vssd1 vccd1 vccd1 _08523_ sky130_fd_sc_hd__a31o_1
XFILLER_36_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17638_ _01915_ vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17569_ rbzero.wall_tracer.rayAddendY\[6\] rbzero.wall_tracer.rayAddendY\[5\] rbzero.wall_tracer.rayAddendY\[4\]
+ rbzero.wall_tracer.rayAddendY\[3\] _01785_ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__o41a_1
X_18981__161 clknet_1_1__leaf__02729_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__inv_2
XFILLER_177_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19308_ rbzero.traced_texa\[-4\] rbzero.texV\[-4\] _02796_ vssd1 vssd1 vccd1 vccd1
+ _02797_ sky130_fd_sc_hd__o21ai_1
XFILLER_143_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19077__247 clknet_1_1__leaf__02739_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__inv_2
XFILLER_173_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20014_ clknet_leaf_92_i_clk _00945_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09825_ rbzero.tex_r1\[17\] rbzero.tex_r1\[18\] _02954_ vssd1 vssd1 vccd1 vccd1 _02961_
+ sky130_fd_sc_hd__mux2_1
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09756_ rbzero.tex_r1\[50\] rbzero.tex_r1\[51\] _02921_ vssd1 vssd1 vccd1 vccd1 _02925_
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10600_ rbzero.map_rom.f2 rbzero.map_rom.f1 rbzero.map_rom.i_col\[4\] vssd1 vssd1
+ vccd1 vccd1 _03396_ sky130_fd_sc_hd__and3_1
XFILLER_70_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11580_ rbzero.tex_b0\[27\] _04155_ _04156_ _03611_ vssd1 vssd1 vccd1 vccd1 _04362_
+ sky130_fd_sc_hd__a31o_1
XFILLER_161_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10531_ rbzero.tex_b0\[4\] rbzero.tex_b0\[3\] _03324_ vssd1 vssd1 vccd1 vccd1 _03333_
+ sky130_fd_sc_hd__mux2_1
XFILLER_161_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13250_ _05469_ _05956_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__nor2_1
X_10462_ rbzero.tex_b0\[37\] rbzero.tex_b0\[36\] _03291_ vssd1 vssd1 vccd1 vccd1 _03297_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19136__300 clknet_1_0__leaf__02745_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__inv_2
XFILLER_171_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12201_ rbzero.wall_tracer.trackDistY\[0\] vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__inv_2
XFILLER_108_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13181_ _05936_ _05937_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__and2_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10393_ rbzero.tex_b1\[5\] rbzero.tex_b1\[6\] _03254_ vssd1 vssd1 vccd1 vccd1 _03261_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12132_ _04892_ _04893_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16940_ _07494_ _08803_ vssd1 vssd1 vccd1 vccd1 _09546_ sky130_fd_sc_hd__or2_1
XFILLER_123_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12063_ _04832_ _03486_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__nor2_1
XFILLER_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11014_ rbzero.row_render.size\[6\] _03774_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__nor2_1
X_16871_ _09269_ _09383_ vssd1 vssd1 vccd1 vccd1 _09478_ sky130_fd_sc_hd__nand2_1
XFILLER_78_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18610_ _02524_ vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15822_ rbzero.traced_texa\[2\] _08461_ _08462_ rbzero.wall_tracer.visualWallDist\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__a22o_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19590_ clknet_leaf_39_i_clk _00521_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18541_ rbzero.pov.spi_buffer\[39\] rbzero.pov.spi_buffer\[40\] _02488_ vssd1 vssd1
+ vccd1 vccd1 _02489_ sky130_fd_sc_hd__mux2_1
XFILLER_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15753_ _08311_ _08434_ _04832_ vssd1 vssd1 vccd1 vccd1 _08436_ sky130_fd_sc_hd__a21o_1
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12965_ _05718_ _05720_ _05721_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__a21o_1
XFILLER_79_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19182__342 clknet_1_0__leaf__02749_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__inv_2
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14704_ _07381_ _07390_ _07391_ vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__a21bo_1
X_11916_ net24 net25 vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__nand2_1
X_15684_ _06997_ _08252_ _08366_ vssd1 vssd1 vccd1 vccd1 _08367_ sky130_fd_sc_hd__or3_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18472_ _02452_ vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _05647_ _05652_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__and2b_1
XFILLER_79_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _07312_ _07320_ _07322_ vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__a21o_1
XFILLER_127_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17423_ _01719_ _01720_ _03486_ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__a21oi_1
XFILLER_54_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11847_ net12 net11 vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__nor2_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14566_ _06873_ _06875_ _07049_ _06857_ vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__o22ai_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _01669_ vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__clkbuf_1
X_11778_ _04552_ _04314_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__nand2_1
XFILLER_186_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16305_ _08910_ _08916_ vssd1 vssd1 vccd1 vccd1 _08917_ sky130_fd_sc_hd__nand2_1
X_13517_ _06237_ _06251_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__nor2_1
X_10729_ gpout0.vpos\[7\] vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__buf_4
X_17285_ _01609_ _01610_ _01611_ vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__a21o_1
XFILLER_201_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14497_ _07157_ vssd1 vssd1 vccd1 vccd1 _07185_ sky130_fd_sc_hd__clkbuf_4
XFILLER_173_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16236_ _08785_ _08764_ vssd1 vssd1 vccd1 vccd1 _08848_ sky130_fd_sc_hd__or2b_1
XFILLER_16_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13448_ _06194_ _06204_ vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16167_ _08777_ _08778_ vssd1 vssd1 vccd1 vccd1 _08780_ sky130_fd_sc_hd__and2_1
XFILLER_142_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13379_ _06119_ _06134_ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__and2_1
XFILLER_86_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15118_ _07372_ _07475_ vssd1 vssd1 vccd1 vccd1 _07806_ sky130_fd_sc_hd__and2b_2
X_16098_ _08427_ _08710_ vssd1 vssd1 vccd1 vccd1 _08712_ sky130_fd_sc_hd__or2_1
XFILLER_88_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19926_ net155 _00857_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[6\] sky130_fd_sc_hd__dfxtp_1
X_15049_ _07734_ _07736_ vssd1 vssd1 vccd1 vccd1 _07737_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_74_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19857_ clknet_leaf_21_i_clk _00788_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_18808_ rbzero.debug_overlay.facingY\[0\] _02634_ vssd1 vssd1 vccd1 vccd1 _02665_
+ sky130_fd_sc_hd__and2_1
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19788_ clknet_leaf_87_i_clk _00719_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[70\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_89_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_110_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18739_ rbzero.debug_overlay.playerY\[3\] _02614_ vssd1 vssd1 vccd1 vccd1 _02619_
+ sky130_fd_sc_hd__or2_1
XFILLER_97_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_12_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_180_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18905__92 clknet_1_1__leaf__02441_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__inv_2
XFILLER_192_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20494_ clknet_leaf_42_i_clk _01425_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19131__296 clknet_1_1__leaf__02744_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__inv_2
X_09808_ rbzero.tex_r1\[25\] rbzero.tex_r1\[26\] _02943_ vssd1 vssd1 vccd1 vccd1 _02952_
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18988__167 clknet_1_0__leaf__02730_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__inv_2
X_09739_ rbzero.tex_r1\[58\] rbzero.tex_r1\[59\] _02910_ vssd1 vssd1 vccd1 vccd1 _02916_
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ _05494_ _05480_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__nand2_1
XFILLER_83_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ rbzero.row_render.texu\[5\] _02899_ _04480_ _03526_ vssd1 vssd1 vccd1 vccd1
+ _04481_ sky130_fd_sc_hd__o211a_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _05372_ _05409_ _05421_ _05437_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__o22a_1
XFILLER_187_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _03492_ rbzero.wall_tracer.stepDistY\[0\] _04949_ vssd1 vssd1 vccd1 vccd1
+ _07108_ sky130_fd_sc_hd__a21oi_1
X_11632_ _04411_ _04412_ _03656_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__mux2_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14351_ _07024_ vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__buf_2
XFILLER_195_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11563_ rbzero.tex_b0\[42\] _03649_ _03823_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__a21o_1
XFILLER_7_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13302_ _06008_ _05988_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__or2_1
XFILLER_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17070_ _09256_ _09229_ vssd1 vssd1 vccd1 vccd1 _09675_ sky130_fd_sc_hd__nor2_1
X_10514_ _02982_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__clkbuf_4
X_14282_ _06966_ vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__clkbuf_4
XFILLER_196_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11494_ rbzero.tex_g1\[53\] rbzero.tex_g1\[52\] _04247_ vssd1 vssd1 vccd1 vccd1 _04277_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16021_ _08633_ _08634_ vssd1 vssd1 vccd1 vccd1 _08635_ sky130_fd_sc_hd__nand2_1
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13233_ _05517_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__clkbuf_4
XFILLER_109_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10445_ rbzero.tex_b0\[45\] rbzero.tex_b0\[44\] _03280_ vssd1 vssd1 vccd1 vccd1 _03288_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13164_ _05870_ _05920_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__or2_1
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10376_ rbzero.tex_b1\[13\] rbzero.tex_b1\[14\] _03243_ vssd1 vssd1 vccd1 vccd1 _03252_
+ sky130_fd_sc_hd__mux2_1
X_12115_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[9\] _04873_
+ _04875_ _04876_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__o221a_1
XFILLER_97_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17972_ rbzero.pov.spi_buffer\[39\] rbzero.pov.ready_buffer\[39\] _02186_ vssd1 vssd1
+ vccd1 vccd1 _02187_ sky130_fd_sc_hd__mux2_1
X_13095_ _05764_ _05800_ _05849_ _05851_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_111_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19711_ clknet_leaf_2_i_clk _00642_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16923_ _09527_ _09462_ _09528_ vssd1 vssd1 vccd1 vccd1 _09529_ sky130_fd_sc_hd__a21oi_2
XFILLER_133_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12046_ _04810_ _04813_ _04818_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__a21o_1
XFILLER_46_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19642_ clknet_leaf_51_i_clk _00573_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16854_ _09345_ _09346_ _09348_ vssd1 vssd1 vccd1 vccd1 _09461_ sky130_fd_sc_hd__o21ai_1
XFILLER_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ rbzero.traced_texa\[-10\] _08457_ _08453_ rbzero.wall_tracer.visualWallDist\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__a22o_1
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19573_ clknet_leaf_41_i_clk _00504_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_16785_ _09391_ _09392_ vssd1 vssd1 vccd1 vccd1 _09393_ sky130_fd_sc_hd__nand2_1
XFILLER_168_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13997_ _05380_ _06699_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__or2_1
XFILLER_19_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18524_ rbzero.pov.spi_buffer\[31\] rbzero.pov.spi_buffer\[32\] _02477_ vssd1 vssd1
+ vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
XFILLER_46_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15736_ _08417_ _08418_ vssd1 vssd1 vccd1 vccd1 _08419_ sky130_fd_sc_hd__nor2_1
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12948_ _05433_ _05536_ vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__nor2_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19108__276 clknet_1_1__leaf__02741_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__inv_2
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18455_ _02442_ vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__clkbuf_4
X_15667_ _08348_ _08349_ vssd1 vssd1 vccd1 vccd1 _08350_ sky130_fd_sc_hd__nor2_1
X_12879_ _05513_ _05634_ _05635_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__or3_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17406_ rbzero.debug_overlay.vplaneY\[-9\] rbzero.wall_tracer.rayAddendY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__nand2_1
XFILLER_61_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14618_ _07300_ _07295_ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__or2b_1
XFILLER_194_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15598_ _08128_ _08156_ _08154_ vssd1 vssd1 vccd1 vccd1 _08282_ sky130_fd_sc_hd__a21oi_2
XFILLER_14_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14549_ _07234_ _07236_ _07233_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__a21boi_1
XFILLER_18_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17337_ rbzero.spi_registers.spi_cmd\[1\] vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__inv_2
XFILLER_105_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17268_ _01598_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__inv_2
XFILLER_88_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16219_ _08721_ _08831_ vssd1 vssd1 vccd1 vccd1 _08832_ sky130_fd_sc_hd__xor2_4
XFILLER_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17199_ _01534_ _01538_ _01539_ _01527_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__a31o_1
XFILLER_115_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19189__348 clknet_1_1__leaf__02750_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__inv_2
X_19909_ clknet_leaf_20_i_clk _00840_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_vshift
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20477_ clknet_leaf_63_i_clk _01408_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10230_ _03175_ vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10161_ rbzero.tex_g0\[52\] rbzero.tex_g0\[51\] _03132_ vssd1 vssd1 vccd1 vccd1 _03139_
+ sky130_fd_sc_hd__mux2_1
XFILLER_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10092_ rbzero.tex_g1\[20\] rbzero.tex_g1\[21\] _03095_ vssd1 vssd1 vccd1 vccd1 _03103_
+ sky130_fd_sc_hd__mux2_1
XFILLER_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13920_ _06097_ _06605_ _05395_ vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__o21ai_2
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13851_ _06474_ _06509_ _06470_ _06557_ vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__a211o_1
XFILLER_74_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12802_ _05505_ _05557_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__nand2_1
XFILLER_74_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16570_ _09178_ _09179_ vssd1 vssd1 vccd1 vccd1 _09180_ sky130_fd_sc_hd__nor2_1
X_13782_ _06531_ _06538_ vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__or2_1
XFILLER_76_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10994_ _03778_ _03779_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__and2_1
XFILLER_16_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15521_ _07235_ _07333_ vssd1 vssd1 vccd1 vccd1 _08205_ sky130_fd_sc_hd__nor2_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _05443_ _05404_ _05425_ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__and3_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15452_ _08131_ _08136_ vssd1 vssd1 vccd1 vccd1 _08137_ sky130_fd_sc_hd__xnor2_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18240_ rbzero.spi_registers.got_new_vshift _02262_ vssd1 vssd1 vccd1 vccd1 _02348_
+ sky130_fd_sc_hd__nand2_2
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _05269_ _05329_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__nand2_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _04947_ rbzero.wall_tracer.stepDistX\[-2\] _07087_ _07090_ vssd1 vssd1 vccd1
+ vccd1 _07091_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_169_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11615_ _04395_ _03998_ _03643_ rbzero.row_render.wall\[1\] vssd1 vssd1 vccd1 vccd1
+ _04396_ sky130_fd_sc_hd__o211a_1
XFILLER_169_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15383_ _07971_ _07989_ _08067_ vssd1 vssd1 vccd1 vccd1 _08068_ sky130_fd_sc_hd__a21bo_1
X_18171_ rbzero.spi_registers.new_mapd\[7\] _02290_ _02303_ _02301_ vssd1 vssd1 vccd1
+ vccd1 _00770_ sky130_fd_sc_hd__o211a_1
X_12595_ _05317_ _05343_ _05346_ _05347_ _05351_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__a221o_1
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17122_ _01463_ _01465_ vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14334_ rbzero.debug_overlay.playerX\[-2\] vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__inv_2
X_11546_ rbzero.tex_b0\[55\] _04155_ _04156_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__and3_1
XFILLER_117_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17053_ _09589_ _09590_ _09592_ vssd1 vssd1 vccd1 vccd1 _09658_ sky130_fd_sc_hd__o21ai_1
XFILLER_184_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14265_ rbzero.wall_tracer.state\[3\] _06682_ _06685_ _06952_ _06859_ vssd1 vssd1
+ vccd1 vccd1 _06953_ sky130_fd_sc_hd__o311a_1
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11477_ _03726_ _04257_ _04258_ _04259_ _03671_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__o221a_1
X_16004_ _08233_ _08359_ vssd1 vssd1 vccd1 vccd1 _08618_ sky130_fd_sc_hd__or2_1
Xclkbuf_0__02742_ _02742_ vssd1 vssd1 vccd1 vccd1 clknet_0__02742_ sky130_fd_sc_hd__clkbuf_16
X_13216_ _05921_ _05951_ _05971_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__and3_1
XFILLER_48_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10428_ rbzero.tex_b0\[53\] rbzero.tex_b0\[52\] _03269_ vssd1 vssd1 vccd1 vccd1 _03279_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14196_ _05096_ _05128_ _05091_ _06883_ vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__and4_1
XFILLER_98_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _05902_ _05903_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__and2b_1
X_10359_ _03072_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__clkbuf_4
XFILLER_135_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13078_ _05767_ _05832_ _05834_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__nor3_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955_ rbzero.pov.spi_buffer\[31\] rbzero.pov.ready_buffer\[31\] _02175_ vssd1 vssd1
+ vccd1 vccd1 _02178_ sky130_fd_sc_hd__mux2_1
XFILLER_140_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16906_ _09511_ _09512_ vssd1 vssd1 vccd1 vccd1 _09513_ sky130_fd_sc_hd__nor2_1
X_12029_ _04798_ _04800_ _04801_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__o21a_1
XFILLER_39_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17886_ rbzero.spi_registers.spi_counter\[6\] _02137_ _02140_ vssd1 vssd1 vccd1 vccd1
+ _00648_ sky130_fd_sc_hd__a21oi_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19625_ clknet_leaf_46_i_clk _00556_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16837_ _09232_ _09337_ _09338_ _09340_ vssd1 vssd1 vccd1 vccd1 _09444_ sky130_fd_sc_hd__a22o_1
XFILLER_76_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19556_ clknet_leaf_10_i_clk _00487_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[6\] sky130_fd_sc_hd__dfxtp_1
X_16768_ _09270_ _09271_ _09273_ vssd1 vssd1 vccd1 vccd1 _09376_ sky130_fd_sc_hd__a21bo_1
XFILLER_81_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18507_ rbzero.pov.spi_buffer\[23\] rbzero.pov.spi_buffer\[24\] _02466_ vssd1 vssd1
+ vccd1 vccd1 _02471_ sky130_fd_sc_hd__mux2_1
XFILLER_62_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15719_ _08400_ _08401_ vssd1 vssd1 vccd1 vccd1 _08402_ sky130_fd_sc_hd__nand2_1
XFILLER_94_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19487_ clknet_leaf_58_i_clk _00433_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-6\]
+ sky130_fd_sc_hd__dfxtp_2
X_16699_ _09304_ _09306_ _09307_ vssd1 vssd1 vccd1 vccd1 _09308_ sky130_fd_sc_hd__a21oi_4
XFILLER_22_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18369_ rbzero.pov.spi_counter\[3\] _02423_ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__nand2_1
XFILLER_187_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20400_ net460 _01331_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20331_ net391 _01262_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20262_ net322 _01193_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20193_ net253 _01124_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02731_ clknet_0__02731_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02731_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ _03702_ _04183_ _03624_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__a21o_1
XFILLER_166_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12380_ _05135_ _05136_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__xnor2_2
XFILLER_197_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_70 net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11331_ _03902_ _03901_ _04097_ _04115_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__o22a_1
XFILLER_158_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14050_ _06784_ vssd1 vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__clkbuf_4
XFILLER_158_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11262_ _04041_ _04043_ _04046_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__o21ai_1
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13001_ _05755_ _05756_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__and2b_1
XFILLER_107_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10213_ rbzero.tex_g0\[28\] rbzero.tex_g0\[27\] _03166_ vssd1 vssd1 vccd1 vccd1 _03167_
+ sky130_fd_sc_hd__mux2_1
XFILLER_106_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11193_ rbzero.tex_r1\[31\] _03936_ _03977_ _03726_ vssd1 vssd1 vccd1 vccd1 _03978_
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10144_ rbzero.tex_g0\[60\] rbzero.tex_g0\[59\] _03050_ vssd1 vssd1 vccd1 vccd1 _03130_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17740_ rbzero.wall_tracer.rayAddendX\[2\] _00013_ _02004_ _02009_ vssd1 vssd1 vccd1
+ vccd1 _00633_ sky130_fd_sc_hd__o22a_1
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10075_ rbzero.tex_g1\[28\] rbzero.tex_g1\[29\] _03084_ vssd1 vssd1 vccd1 vccd1 _03094_
+ sky130_fd_sc_hd__mux2_1
X_14952_ _07636_ _07638_ _07639_ vssd1 vssd1 vccd1 vccd1 _07640_ sky130_fd_sc_hd__a21oi_1
XFILLER_43_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13903_ _05265_ _05271_ _06652_ _06657_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__a31o_1
X_17671_ _01942_ _01943_ _01945_ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__o21ai_1
XFILLER_47_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14883_ _07529_ _07570_ vssd1 vssd1 vccd1 vccd1 _07571_ sky130_fd_sc_hd__or2_1
XFILLER_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19410_ rbzero.debug_overlay.vplaneY\[-9\] rbzero.wall_tracer.rayAddendY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__or2_1
XFILLER_63_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16622_ _07333_ vssd1 vssd1 vccd1 vccd1 _09231_ sky130_fd_sc_hd__buf_2
X_13834_ _06577_ _06590_ _06578_ _06218_ vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19341_ _02822_ _02823_ _02824_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__and3_1
X_16553_ _09161_ _09162_ vssd1 vssd1 vccd1 vccd1 _09163_ sky130_fd_sc_hd__and2_1
X_13765_ _06487_ _06519_ _06521_ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__a21bo_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10977_ _03688_ _03754_ _03762_ _03718_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__a31o_1
XFILLER_31_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15504_ _08087_ _08089_ _08090_ _08074_ vssd1 vssd1 vccd1 vccd1 _08188_ sky130_fd_sc_hd__a2bb2o_1
X_12716_ _05443_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__buf_2
XFILLER_43_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19272_ _02764_ _02765_ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__and2_1
X_16484_ _08983_ _08984_ _08981_ vssd1 vssd1 vccd1 vccd1 _09094_ sky130_fd_sc_hd__a21oi_1
X_13696_ _06122_ _06070_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__nor2_1
XFILLER_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18223_ _02334_ _02336_ vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__and2_1
XFILLER_175_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15435_ _07997_ _08118_ _08119_ vssd1 vssd1 vccd1 vccd1 _08120_ sky130_fd_sc_hd__o21a_1
X_12647_ _05369_ _05399_ _05401_ _05403_ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__o31a_4
XFILLER_31_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15366_ _08048_ _08051_ vssd1 vssd1 vccd1 vccd1 _08052_ sky130_fd_sc_hd__xnor2_4
X_18154_ rbzero.spi_registers.new_mapd\[11\] _02290_ _02294_ _02275_ vssd1 vssd1 vccd1
+ vccd1 _00762_ sky130_fd_sc_hd__o211a_1
X_12578_ _05210_ _05334_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__nor2_1
XFILLER_200_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17105_ rbzero.wall_tracer.trackDistX\[9\] rbzero.wall_tracer.stepDistX\[9\] vssd1
+ vssd1 vccd1 vccd1 _09710_ sky130_fd_sc_hd__nand2_1
XFILLER_157_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14317_ _04839_ rbzero.wall_tracer.stepDistX\[-8\] _07001_ _07004_ vssd1 vssd1 vccd1
+ vccd1 _07005_ sky130_fd_sc_hd__a2bb2o_4
X_11529_ _03848_ _04018_ _04310_ _04311_ _03897_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__a41o_1
XFILLER_116_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15297_ _07981_ _07982_ vssd1 vssd1 vccd1 vccd1 _07983_ sky130_fd_sc_hd__xnor2_1
X_18085_ _02247_ vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__clkbuf_1
XFILLER_116_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17036_ _09639_ _09640_ vssd1 vssd1 vccd1 vccd1 _09641_ sky130_fd_sc_hd__xor2_2
X_14248_ rbzero.wall_tracer.state\[3\] _06935_ vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__nand2_1
Xclkbuf_0__02725_ _02725_ vssd1 vssd1 vccd1 vccd1 clknet_0__02725_ sky130_fd_sc_hd__clkbuf_16
XFILLER_125_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14179_ _03491_ rbzero.wall_tracer.stepDistY\[-10\] _04948_ vssd1 vssd1 vccd1 vccd1
+ _06867_ sky130_fd_sc_hd__a21oi_1
XFILLER_113_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ clknet_1_1__leaf__02440_ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__buf_1
XFILLER_61_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ rbzero.pov.spi_buffer\[23\] rbzero.pov.ready_buffer\[23\] _02164_ vssd1 vssd1
+ vccd1 vccd1 _02169_ sky130_fd_sc_hd__mux2_1
XFILLER_78_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17869_ rbzero.spi_registers.spi_counter\[2\] _02102_ vssd1 vssd1 vccd1 vccd1 _02128_
+ sky130_fd_sc_hd__or2_1
XFILLER_93_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19608_ clknet_leaf_54_i_clk _00539_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_199_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19539_ clknet_leaf_58_i_clk _00010_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20314_ net374 _01245_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20245_ net305 _01176_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09987_ _03047_ vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__clkbuf_1
X_20176_ net236 _01107_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10900_ _03648_ _03658_ _03672_ _03680_ _03685_ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__o221a_1
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11880_ _04507_ _04508_ _03520_ _03515_ _04612_ net11 vssd1 vssd1 vccd1 vccd1 _04656_
+ sky130_fd_sc_hd__mux4_1
Xtop_ew_algofoogle_109 vssd1 vssd1 vccd1 vccd1 ones[2] top_ew_algofoogle_109/LO sky130_fd_sc_hd__conb_1
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10831_ _03616_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__clkbuf_8
XFILLER_26_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13550_ _06304_ _06306_ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__nor2_1
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10762_ rbzero.traced_texVinit\[3\] rbzero.spi_registers.vshift\[0\] vssd1 vssd1
+ vccd1 vccd1 _03548_ sky130_fd_sc_hd__nand2_1
XFILLER_52_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12501_ _05094_ _05227_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__xnor2_2
XFILLER_201_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13481_ _05301_ _05527_ _06055_ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__or3_1
XFILLER_201_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10693_ _03484_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__buf_6
XFILLER_200_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15220_ _07760_ _07762_ vssd1 vssd1 vccd1 vccd1 _07907_ sky130_fd_sc_hd__nor2_1
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12432_ _05186_ _05188_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__xor2_2
XFILLER_40_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15151_ _07836_ _07837_ vssd1 vssd1 vccd1 vccd1 _07838_ sky130_fd_sc_hd__nand2_1
X_12363_ _03487_ _05107_ _05109_ _05114_ _05119_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__a2111o_4
XFILLER_138_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14102_ rbzero.wall_tracer.visualWallDist\[10\] _03496_ _06815_ _03498_ vssd1 vssd1
+ vccd1 vccd1 _00449_ sky130_fd_sc_hd__o211a_1
XFILLER_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11314_ rbzero.debug_overlay.vplaneX\[-1\] _04093_ _04056_ rbzero.debug_overlay.vplaneX\[-2\]
+ _04098_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__a221o_1
X_15082_ _07764_ _07769_ vssd1 vssd1 vccd1 vccd1 _07770_ sky130_fd_sc_hd__xor2_2
XFILLER_180_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12294_ _05034_ _05037_ _05046_ _05048_ _05050_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__a311o_1
XFILLER_154_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18910_ clknet_1_0__leaf__02440_ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__buf_1
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14033_ _06771_ vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__inv_2
X_11245_ _04005_ _04029_ _03848_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__o21a_1
XFILLER_180_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19890_ clknet_leaf_20_i_clk _00821_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_106_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18841_ rbzero.debug_overlay.vplaneY\[-7\] _02660_ vssd1 vssd1 vccd1 vccd1 _02683_
+ sky130_fd_sc_hd__or2_1
X_11176_ rbzero.tex_r1\[5\] _03919_ _03926_ _03673_ vssd1 vssd1 vccd1 vccd1 _03961_
+ sky130_fd_sc_hd__a31o_1
XFILLER_132_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__02441_ _02441_ vssd1 vssd1 vccd1 vccd1 clknet_0__02441_ sky130_fd_sc_hd__clkbuf_16
X_10127_ _03121_ vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__clkbuf_1
X_18772_ _02633_ vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__buf_2
XFILLER_110_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15984_ _07011_ _08318_ _08317_ _08597_ vssd1 vssd1 vccd1 vccd1 _08598_ sky130_fd_sc_hd__a31o_1
XFILLER_0_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17723_ _01992_ _01993_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__nor2_1
X_14935_ _07049_ _07213_ vssd1 vssd1 vccd1 vccd1 _07623_ sky130_fd_sc_hd__or2_1
X_10058_ _03085_ vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17654_ rbzero.debug_overlay.vplaneX\[-9\] _01930_ _03484_ vssd1 vssd1 vccd1 vccd1
+ _01931_ sky130_fd_sc_hd__mux2_1
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14866_ _06939_ _06954_ _07156_ _07177_ vssd1 vssd1 vccd1 vccd1 _07554_ sky130_fd_sc_hd__nor4_1
XFILLER_90_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16605_ _08107_ _08191_ vssd1 vssd1 vccd1 vccd1 _09214_ sky130_fd_sc_hd__nor2_1
XFILLER_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13817_ _06573_ _06568_ _06227_ vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__a21o_1
X_17585_ _01757_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__inv_2
XFILLER_32_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14797_ _07482_ _07483_ _07484_ vssd1 vssd1 vccd1 vccd1 _07485_ sky130_fd_sc_hd__o21ai_1
X_19324_ _02807_ _02808_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__nor2_1
XFILLER_188_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16536_ _09144_ _09145_ vssd1 vssd1 vccd1 vccd1 _09146_ sky130_fd_sc_hd__nor2_1
XFILLER_73_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13748_ _06497_ _06504_ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__nand2_1
XFILLER_32_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16467_ _08952_ _08953_ vssd1 vssd1 vccd1 vccd1 _09078_ sky130_fd_sc_hd__nor2_1
X_13679_ _06397_ _06423_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__xor2_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18206_ _02323_ _02324_ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__and2_1
XFILLER_176_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15418_ _07039_ _07273_ _07141_ _07092_ vssd1 vssd1 vccd1 vccd1 _08103_ sky130_fd_sc_hd__or4_1
XFILLER_192_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16398_ _06858_ vssd1 vssd1 vccd1 vccd1 _09009_ sky130_fd_sc_hd__buf_2
XFILLER_185_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18137_ _02279_ _02259_ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__and2_1
X_15349_ _08032_ _08034_ vssd1 vssd1 vccd1 vccd1 _08035_ sky130_fd_sc_hd__xor2_2
XFILLER_117_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18068_ rbzero.spi_registers.spi_buffer\[10\] rbzero.spi_registers.spi_buffer\[9\]
+ _02226_ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__mux2_1
XFILLER_176_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09910_ _03007_ vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__clkbuf_1
X_17019_ _09521_ _09524_ _09522_ vssd1 vssd1 vccd1 vccd1 _09625_ sky130_fd_sc_hd__o21ai_1
XFILLER_171_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09841_ _02969_ vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__clkbuf_1
X_20030_ clknet_leaf_85_i_clk _00961_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09772_ _02933_ vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__clkbuf_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11030_ _03460_ _03803_ _03801_ _03466_ _03815_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__a221o_1
X_20228_ net288 _01159_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20159_ net219 _01090_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12981_ _05493_ _05535_ _05737_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__or3b_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ _07393_ _07406_ _07407_ vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__a21boi_2
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11932_ _04672_ net67 _04706_ net25 vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__a211o_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ net124 _04626_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__nand2_2
X_14651_ _07329_ _07338_ vssd1 vssd1 vccd1 vccd1 _07339_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10814_ _03572_ _03575_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__nand2_1
X_13602_ _06343_ _06350_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__xor2_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _01677_ vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__clkbuf_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14582_ _07257_ vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__buf_2
X_11794_ net20 net19 vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__nor2_1
XFILLER_186_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16321_ _08808_ _08810_ vssd1 vssd1 vccd1 vccd1 _08933_ sky130_fd_sc_hd__and2b_1
XFILLER_159_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13533_ _05862_ _05988_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__nor2_1
X_10745_ gpout0.vpos\[7\] gpout0.vpos\[6\] _03519_ vssd1 vssd1 vccd1 vccd1 _03531_
+ sky130_fd_sc_hd__or3_1
XFILLER_186_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16252_ _07993_ _07857_ _08769_ _08863_ vssd1 vssd1 vccd1 vccd1 _08864_ sky130_fd_sc_hd__o31ai_1
XFILLER_146_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13464_ _06194_ _06204_ _06220_ vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__a21oi_1
X_10676_ _03459_ _03468_ _03470_ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__a21o_1
XFILLER_199_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15203_ _07888_ _07889_ vssd1 vssd1 vccd1 vccd1 _07890_ sky130_fd_sc_hd__nand2_1
X_12415_ _03489_ _05171_ _05170_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__a21oi_1
X_16183_ _08794_ _08795_ vssd1 vssd1 vccd1 vccd1 _08796_ sky130_fd_sc_hd__and2_1
XFILLER_138_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13395_ _06008_ _05995_ _06151_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__or3b_1
XFILLER_154_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12346_ _03479_ _04894_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__nand2_1
X_15134_ _07812_ _07821_ vssd1 vssd1 vccd1 vccd1 _07822_ sky130_fd_sc_hd__or2_1
X_19942_ net171 _00873_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15065_ _03492_ rbzero.wall_tracer.stepDistY\[5\] _04948_ vssd1 vssd1 vccd1 vccd1
+ _07753_ sky130_fd_sc_hd__a21oi_1
XFILLER_181_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12277_ _05032_ _05033_ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__nor2_1
XFILLER_5_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14016_ _06630_ _06757_ vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__or2_1
X_11228_ _03852_ _03782_ _04008_ _04012_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__a31o_1
X_19873_ clknet_leaf_22_i_clk _00804_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18824_ _04102_ _02634_ vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__and2_1
XFILLER_110_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11159_ rbzero.tex_r1\[42\] _03620_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__or2_1
XFILLER_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18755_ rbzero.pov.ready _02607_ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__and2_1
XFILLER_48_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15967_ _08562_ _08581_ _08582_ _08522_ vssd1 vssd1 vccd1 vccd1 _08583_ sky130_fd_sc_hd__a31o_1
XFILLER_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17706_ _04102_ rbzero.debug_overlay.vplaneX\[-8\] vssd1 vssd1 vccd1 vccd1 _01978_
+ sky130_fd_sc_hd__nand2_1
X_14918_ _07584_ _07604_ vssd1 vssd1 vccd1 vccd1 _07606_ sky130_fd_sc_hd__nand2_1
XFILLER_76_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18686_ rbzero.debug_overlay.playerX\[5\] rbzero.debug_overlay.playerX\[4\] _02570_
+ _02540_ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__o31ai_1
X_15898_ _08487_ vssd1 vssd1 vccd1 vccd1 _08522_ sky130_fd_sc_hd__clkbuf_4
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17637_ _01914_ rbzero.wall_tracer.mapY\[5\] _05006_ vssd1 vssd1 vccd1 vccd1 _01915_
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14849_ _07491_ _07490_ vssd1 vssd1 vccd1 vccd1 _07537_ sky130_fd_sc_hd__nand2_1
XFILLER_1_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17568_ _01829_ _01830_ _01842_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__nor3_1
XFILLER_189_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19307_ rbzero.traced_texa\[-4\] rbzero.texV\[-4\] _02792_ vssd1 vssd1 vccd1 vccd1
+ _02796_ sky130_fd_sc_hd__a21o_1
X_16519_ _09127_ _09128_ vssd1 vssd1 vccd1 vccd1 _09129_ sky130_fd_sc_hd__nand2_1
XFILLER_108_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17499_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.debug_overlay.vplaneY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__nor2_1
XFILLER_143_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20013_ clknet_leaf_92_i_clk _00944_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09824_ _02960_ vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09755_ _02924_ vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10530_ _03332_ vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10461_ _03296_ vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12200_ rbzero.wall_tracer.trackDistY\[2\] vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__inv_2
XFILLER_159_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13180_ _05873_ _05911_ _05935_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__nand3_1
XFILLER_109_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10392_ _03260_ vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12131_ _04858_ _04862_ _04863_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__a21oi_1
XFILLER_135_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12062_ _04831_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__buf_4
XFILLER_96_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19246__20 clknet_1_0__leaf__02755_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__inv_2
XFILLER_81_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11013_ _02900_ _03798_ _03797_ _02902_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__a22o_1
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16870_ _09361_ _09370_ _09368_ vssd1 vssd1 vccd1 vccd1 _09477_ sky130_fd_sc_hd__a21o_1
XFILLER_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15821_ rbzero.traced_texa\[1\] _08461_ _08462_ rbzero.wall_tracer.visualWallDist\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__a22o_1
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18540_ _02443_ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__clkbuf_4
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _08311_ _08434_ vssd1 vssd1 vccd1 vccd1 _08435_ sky130_fd_sc_hd__nor2_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _05716_ _05717_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__nor2_1
XFILLER_92_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ _07389_ _07383_ vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__or2b_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18471_ rbzero.pov.spi_buffer\[6\] rbzero.pov.spi_buffer\[7\] _02444_ vssd1 vssd1
+ vccd1 vccd1 _02452_ sky130_fd_sc_hd__mux2_1
X_11915_ _04682_ _04684_ _04689_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__a21oi_2
X_15683_ _07494_ _07198_ vssd1 vssd1 vccd1 vccd1 _08366_ sky130_fd_sc_hd__or2_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _05493_ _05551_ _05648_ _05650_ _05651_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__o32ai_4
XFILLER_33_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _01716_ _01717_ _01718_ vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__o21ai_1
X_14634_ _07261_ _07321_ vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__nand2_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11846_ net10 net9 vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__nor2_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ rbzero.spi_registers.new_mapd\[5\] rbzero.spi_registers.spi_buffer\[5\] _01663_
+ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__mux2_1
X_14565_ _06874_ _07013_ _07049_ vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__or3_1
X_11777_ _04552_ net67 _04553_ net19 vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__a211o_1
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _08914_ _08915_ vssd1 vssd1 vccd1 vccd1 _08916_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13516_ _06229_ _06272_ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__xnor2_1
X_10728_ gpout0.hpos\[8\] _03513_ gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 _03514_
+ sky130_fd_sc_hd__a21oi_2
X_17284_ _01612_ vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__inv_2
X_14496_ _07154_ _07157_ _07179_ _07183_ _07168_ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__o32a_1
XFILLER_174_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16235_ _08741_ _08758_ _08756_ vssd1 vssd1 vccd1 vccd1 _08847_ sky130_fd_sc_hd__a21o_1
XFILLER_146_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13447_ _06202_ _06203_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__xor2_1
X_10659_ _03432_ _03445_ _03454_ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__o21ba_1
XFILLER_173_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19002__180 clknet_1_1__leaf__02731_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__inv_2
XFILLER_103_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16166_ _08777_ _08778_ vssd1 vssd1 vccd1 vccd1 _08779_ sky130_fd_sc_hd__nor2_1
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13378_ _06119_ _06134_ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__nor2_1
XFILLER_126_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15117_ _07803_ _07804_ vssd1 vssd1 vccd1 vccd1 _07805_ sky130_fd_sc_hd__xor2_4
X_12329_ _05082_ _05085_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__xnor2_2
XFILLER_114_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16097_ _08427_ _08710_ vssd1 vssd1 vccd1 vccd1 _08711_ sky130_fd_sc_hd__nand2_1
XFILLER_114_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15048_ _07735_ _06993_ vssd1 vssd1 vccd1 vccd1 _07736_ sky130_fd_sc_hd__nor2_1
X_19925_ net154 _00856_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[5\] sky130_fd_sc_hd__dfxtp_1
X_19856_ clknet_leaf_23_i_clk _00787_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18807_ rbzero.pov.ready_buffer\[30\] _02663_ _02664_ _02643_ vssd1 vssd1 vccd1 vccd1
+ _01045_ sky130_fd_sc_hd__o211a_1
XFILLER_95_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19787_ clknet_leaf_86_i_clk _00718_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[69\]
+ sky130_fd_sc_hd__dfxtp_1
X_16999_ _09531_ _09603_ vssd1 vssd1 vccd1 vccd1 _09605_ sky130_fd_sc_hd__or2_1
X_18445__84 clknet_1_0__leaf__02439_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__inv_2
XFILLER_62_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18738_ _03347_ _02587_ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__nor2_1
XFILLER_48_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18669_ rbzero.debug_overlay.playerX\[1\] _02533_ _02565_ _02559_ vssd1 vssd1 vccd1
+ vccd1 _01006_ sky130_fd_sc_hd__a211o_1
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20493_ clknet_leaf_43_i_clk _01424_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09807_ _02951_ vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19166__327 clknet_1_0__leaf__02748_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__inv_2
X_09738_ _02915_ vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11700_ rbzero.row_render.texu\[4\] _02899_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__or2b_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _05294_ _05313_ _05406_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__o21ai_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11631_ rbzero.tex_b1\[35\] rbzero.tex_b1\[34\] _03616_ vssd1 vssd1 vccd1 vccd1 _04412_
+ sky130_fd_sc_hd__mux2_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11562_ rbzero.tex_b0\[43\] _03696_ _03697_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__and3_1
X_14350_ _07005_ _07037_ vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__or2_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10513_ _03323_ vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13301_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14281_ _06954_ vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__buf_4
X_11493_ _04274_ _04275_ _03612_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__mux2_1
XFILLER_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16020_ _08605_ _08606_ _08632_ vssd1 vssd1 vccd1 vccd1 _08634_ sky130_fd_sc_hd__nand3_1
X_13232_ _05472_ _05988_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__or2_1
XFILLER_196_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10444_ _03287_ vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13163_ _05861_ _05919_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__xnor2_1
X_10375_ _03251_ vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12114_ rbzero.debug_overlay.facingY\[0\] rbzero.wall_tracer.rayAddendY\[8\] vssd1
+ vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__or2_1
XFILLER_2_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13094_ _05765_ _05850_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__xnor2_1
X_17971_ _02142_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__clkbuf_4
XFILLER_124_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19710_ clknet_leaf_72_i_clk _00641_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_16922_ _09437_ _09438_ _09441_ vssd1 vssd1 vccd1 vccd1 _09528_ sky130_fd_sc_hd__o21a_1
X_12045_ _04815_ _04817_ net37 vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__a21bo_1
XFILLER_2_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19641_ clknet_leaf_51_i_clk _00572_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16853_ _09432_ _09459_ vssd1 vssd1 vccd1 vccd1 _09460_ sky130_fd_sc_hd__xor2_1
XFILLER_120_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15804_ rbzero.traced_texa\[-11\] _08457_ _08453_ _06787_ vssd1 vssd1 vccd1 vccd1
+ _00509_ sky130_fd_sc_hd__a22o_1
X_19572_ clknet_leaf_41_i_clk _00503_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_16784_ _09375_ _09390_ vssd1 vssd1 vccd1 vccd1 _09392_ sky130_fd_sc_hd__or2_1
XFILLER_81_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13996_ _06675_ _06684_ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__and2_1
XFILLER_93_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18523_ _02479_ vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__clkbuf_1
X_15735_ _08356_ _08284_ _08416_ vssd1 vssd1 vccd1 vccd1 _08418_ sky130_fd_sc_hd__and3_1
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ _05526_ _05493_ _05535_ _05465_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__or4b_1
XFILLER_34_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18454_ _02415_ _02414_ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__nand2_1
X_15666_ _08346_ _08347_ vssd1 vssd1 vccd1 vccd1 _08349_ sky130_fd_sc_hd__and2_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12878_ _05484_ _05471_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__nor2_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17405_ rbzero.debug_overlay.vplaneY\[-7\] rbzero.wall_tracer.rayAddendY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__nor2_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14617_ _07303_ _07304_ vssd1 vssd1 vccd1 vccd1 _07305_ sky130_fd_sc_hd__xnor2_1
X_11829_ _04507_ _04508_ _03520_ _03515_ _04552_ net17 vssd1 vssd1 vccd1 vccd1 _04606_
+ sky130_fd_sc_hd__mux4_1
X_15597_ _08258_ _08280_ vssd1 vssd1 vccd1 vccd1 _08281_ sky130_fd_sc_hd__xnor2_2
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17336_ _01657_ _01514_ rbzero.wall_tracer.trackDistY\[10\] _01523_ vssd1 vssd1 vccd1
+ vccd1 _00581_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14548_ _07235_ _06993_ vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__nor2_1
XFILLER_14_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17267_ _01595_ _01596_ _01597_ vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__and3_1
XFILLER_174_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14479_ _06860_ _07159_ _07162_ _07166_ _04840_ vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__o221a_1
XFILLER_162_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16218_ _08829_ _08830_ vssd1 vssd1 vccd1 vccd1 _08831_ sky130_fd_sc_hd__nand2_2
XFILLER_128_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17198_ _01536_ _01537_ _01535_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__o21ai_1
X_16149_ _08760_ _08761_ vssd1 vssd1 vccd1 vccd1 _08762_ sky130_fd_sc_hd__nand2_1
XFILLER_103_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19908_ clknet_leaf_19_i_clk _00839_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19839_ clknet_leaf_15_i_clk _00770_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19240__15 clknet_1_0__leaf__02754_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__inv_2
XFILLER_71_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20476_ clknet_leaf_37_i_clk _01407_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10160_ _03138_ vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10091_ _03102_ vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__clkbuf_1
X_18409__51 clknet_1_0__leaf__02436_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__inv_2
XFILLER_0_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13850_ _05271_ _06604_ _06606_ _05356_ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__a211o_1
XFILLER_75_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18424__65 clknet_1_0__leaf__02437_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__inv_2
XFILLER_63_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12801_ _05404_ _05557_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__or2_1
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13781_ _06533_ _06535_ _06537_ vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__o21a_1
XFILLER_56_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10993_ rbzero.row_render.size\[8\] rbzero.row_render.size\[7\] rbzero.row_render.size\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__nand3_1
XFILLER_167_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15520_ _07972_ _07787_ vssd1 vssd1 vccd1 vccd1 _08204_ sky130_fd_sc_hd__nor2_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12732_ _05443_ _05425_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__nor2_4
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15451_ _08132_ _08135_ vssd1 vssd1 vccd1 vccd1 _08136_ sky130_fd_sc_hd__nand2_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _05418_ _05419_ _05270_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_73_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14402_ rbzero.wall_tracer.state\[3\] _06717_ _07089_ _06859_ vssd1 vssd1 vccd1 vccd1
+ _07090_ sky130_fd_sc_hd__o211a_1
XFILLER_187_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11614_ _04198_ _03661_ _03630_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__a21oi_1
X_18170_ rbzero.map_overlay.i_mapdy\[3\] _02292_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__or2_1
X_15382_ _07990_ _07969_ vssd1 vssd1 vccd1 vccd1 _08067_ sky130_fd_sc_hd__or2b_1
XFILLER_168_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12594_ _05348_ _05350_ _05325_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__mux2_1
XFILLER_196_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17121_ _09636_ _01464_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__xor2_1
X_14333_ rbzero.debug_overlay.playerX\[-2\] _06987_ vssd1 vssd1 vccd1 vccd1 _07021_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_195_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11545_ rbzero.tex_b0\[53\] rbzero.tex_b0\[52\] _03732_ vssd1 vssd1 vccd1 vccd1 _04327_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17052_ _09632_ _09656_ vssd1 vssd1 vccd1 vccd1 _09657_ sky130_fd_sc_hd__xnor2_1
XFILLER_144_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11476_ rbzero.tex_g1\[15\] _03729_ _03730_ _03612_ vssd1 vssd1 vccd1 vccd1 _04259_
+ sky130_fd_sc_hd__a31o_1
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14264_ _06849_ _05102_ _06951_ _04830_ vssd1 vssd1 vccd1 vccd1 _06952_ sky130_fd_sc_hd__a211o_1
XFILLER_109_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_88_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16003_ _08227_ _08616_ _08340_ _08206_ vssd1 vssd1 vccd1 vccd1 _08617_ sky130_fd_sc_hd__a22o_1
XFILLER_125_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10427_ _03278_ vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__02741_ _02741_ vssd1 vssd1 vccd1 vccd1 clknet_0__02741_ sky130_fd_sc_hd__clkbuf_16
XFILLER_125_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13215_ _05921_ _05951_ _05971_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__a21oi_1
X_14195_ _05124_ _05102_ _06882_ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__nor3_1
XFILLER_48_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10358_ _03242_ vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__clkbuf_1
X_13146_ _05849_ _05851_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__xor2_2
XFILLER_48_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_11_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13077_ _05797_ _05833_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__nand2_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17954_ _02177_ vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10289_ _03206_ vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__clkbuf_1
X_19114__281 clknet_1_0__leaf__02742_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__inv_2
XFILLER_78_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16905_ _09508_ _09510_ vssd1 vssd1 vccd1 vccd1 _09512_ sky130_fd_sc_hd__and2_1
X_12028_ net35 vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__inv_2
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17885_ rbzero.spi_registers.spi_counter\[6\] _02137_ _02103_ vssd1 vssd1 vccd1 vccd1
+ _02140_ sky130_fd_sc_hd__o21ai_1
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16836_ _09441_ _09442_ vssd1 vssd1 vccd1 vccd1 _09443_ sky130_fd_sc_hd__and2_1
XFILLER_38_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19624_ clknet_leaf_46_i_clk _00555_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_26_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_19_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19555_ clknet_leaf_10_i_clk _00486_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[5\] sky130_fd_sc_hd__dfxtp_1
X_16767_ _09355_ _09374_ vssd1 vssd1 vccd1 vccd1 _09375_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13979_ _05414_ _06720_ _06725_ vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__a21o_2
X_18506_ _02470_ vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15718_ _07175_ _04950_ _03493_ _08399_ _08315_ vssd1 vssd1 vccd1 vccd1 _08401_ sky130_fd_sc_hd__o41ai_1
XFILLER_20_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19486_ clknet_leaf_59_i_clk _00432_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-7\]
+ sky130_fd_sc_hd__dfxtp_2
X_16698_ _09304_ _09306_ _08485_ vssd1 vssd1 vccd1 vccd1 _09307_ sky130_fd_sc_hd__o21ai_1
XFILLER_34_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18437_ clknet_1_0__leaf__02433_ vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__buf_1
X_15649_ _08330_ _08331_ vssd1 vssd1 vccd1 vccd1 _08332_ sky130_fd_sc_hd__nand2_1
XFILLER_181_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18368_ _02423_ _02424_ vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__nor2_1
XFILLER_175_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17319_ _01640_ _01641_ _01642_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__a21oi_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18299_ rbzero.spi_registers.spi_buffer\[3\] rbzero.spi_registers.new_leak\[3\] _02379_
+ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__mux2_1
XFILLER_119_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20330_ net390 _01261_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20261_ net321 _01192_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20192_ net252 _01123_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__02730_ clknet_0__02730_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02730_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_60 _07151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_71 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11330_ _03903_ _04106_ _04114_ _03900_ _03852_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__o32a_1
XFILLER_193_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11261_ gpout0.hpos\[5\] _03466_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__nand2_1
XFILLER_107_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20459_ net139 _01390_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10212_ _03143_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__clkbuf_4
X_13000_ _05755_ _05756_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__xnor2_1
XFILLER_107_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11192_ rbzero.tex_r1\[30\] _03926_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__or2_1
XFILLER_79_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10143_ _03129_ vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10074_ _03093_ vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__clkbuf_1
X_14951_ _07583_ _07607_ vssd1 vssd1 vccd1 vccd1 _07639_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13902_ _06654_ _06656_ _06630_ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__a21o_1
X_17670_ _04102_ rbzero.wall_tracer.rayAddendX\[-4\] _01944_ vssd1 vssd1 vccd1 vccd1
+ _01945_ sky130_fd_sc_hd__o21ai_1
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14882_ _07544_ _07568_ _07569_ vssd1 vssd1 vccd1 vccd1 _07570_ sky130_fd_sc_hd__a21boi_2
XFILLER_48_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16621_ _08862_ _09229_ vssd1 vssd1 vccd1 vccd1 _09230_ sky130_fd_sc_hd__nor2_1
XFILLER_29_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13833_ _06081_ _06196_ _06576_ vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__or3_1
XFILLER_29_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19340_ _02817_ _02820_ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__nand2_1
X_16552_ _09048_ _09155_ _09160_ vssd1 vssd1 vccd1 vccd1 _09162_ sky130_fd_sc_hd__nand3_1
X_13764_ _05805_ _06071_ _06520_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__or3b_1
XFILLER_90_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _03689_ _03757_ _03761_ _03704_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__a211o_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15503_ _08068_ _08091_ _08186_ vssd1 vssd1 vccd1 vccd1 _08187_ sky130_fd_sc_hd__a21bo_1
X_12715_ _05471_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__buf_2
XFILLER_31_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19271_ _02759_ _02765_ _02766_ _02762_ rbzero.texV\[-10\] vssd1 vssd1 vccd1 vccd1
+ _01407_ sky130_fd_sc_hd__a32o_1
X_16483_ _09004_ _08973_ vssd1 vssd1 vccd1 vccd1 _09093_ sky130_fd_sc_hd__or2b_1
XFILLER_16_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13695_ _06409_ _06411_ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18222_ rbzero.color_floor\[0\] rbzero.spi_registers.new_floor\[0\] _02335_ vssd1
+ vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__mux2_1
XFILLER_176_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15434_ _06968_ _06970_ _07137_ _07198_ vssd1 vssd1 vccd1 vccd1 _08119_ sky130_fd_sc_hd__or4_1
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12646_ _05209_ _05376_ _05322_ _05402_ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__or4_1
XFILLER_169_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18153_ rbzero.map_overlay.i_mapdx\[1\] _02292_ vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__or2_1
XFILLER_200_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15365_ _07832_ _08049_ _08050_ _07830_ vssd1 vssd1 vccd1 vccd1 _08051_ sky130_fd_sc_hd__o22a_2
XFILLER_178_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12577_ _05333_ _05300_ _05278_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__a21bo_2
XFILLER_184_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17104_ _09706_ _09707_ _09708_ vssd1 vssd1 vccd1 vccd1 _09709_ sky130_fd_sc_hd__o21ai_2
XFILLER_190_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ _06852_ _06669_ _07003_ _06985_ vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__o211ai_1
XFILLER_129_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18084_ _02107_ rbzero.spi_registers.spi_cmd\[1\] _02245_ vssd1 vssd1 vccd1 vccd1
+ _02247_ sky130_fd_sc_hd__mux2_1
X_11528_ _03860_ _04005_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__nor2_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15296_ _07097_ _07052_ vssd1 vssd1 vccd1 vccd1 _07982_ sky130_fd_sc_hd__or2_1
XFILLER_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17035_ _08889_ _09039_ vssd1 vssd1 vccd1 vccd1 _09640_ sky130_fd_sc_hd__nor2_1
X_14247_ _04901_ _05128_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _06935_ sky130_fd_sc_hd__mux2_1
X_11459_ _04240_ _04241_ _03612_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__02724_ _02724_ vssd1 vssd1 vccd1 vccd1 clknet_0__02724_ sky130_fd_sc_hd__clkbuf_16
XFILLER_131_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14178_ _06865_ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__buf_4
XFILLER_125_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _05636_ _05885_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__xor2_1
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17937_ _02168_ vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17868_ rbzero.spi_registers.spi_counter\[2\] _02112_ _02126_ vssd1 vssd1 vccd1 vccd1
+ _02127_ sky130_fd_sc_hd__a21oi_1
XFILLER_54_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19607_ clknet_leaf_54_i_clk _00538_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
X_16819_ _09351_ _09424_ _09425_ vssd1 vssd1 vccd1 vccd1 _09426_ sky130_fd_sc_hd__a21oi_1
XFILLER_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17799_ _02039_ _02037_ _02050_ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__nor3b_1
XFILLER_54_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18403__46 clknet_1_0__leaf__02435_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__inv_2
XFILLER_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19538_ clknet_leaf_67_i_clk _00009_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_185_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19469_ clknet_leaf_52_i_clk _00415_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20313_ net373 _01244_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20244_ net304 _01175_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20175_ net235 _01106_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09986_ rbzero.tex_r0\[7\] rbzero.tex_r0\[6\] _03039_ vssd1 vssd1 vccd1 vccd1 _03047_
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10830_ _03615_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__buf_6
XFILLER_60_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10761_ rbzero.traced_texVinit\[3\] rbzero.spi_registers.vshift\[0\] vssd1 vssd1
+ vccd1 vccd1 _03547_ sky130_fd_sc_hd__or2_1
XFILLER_201_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12500_ _05202_ _05203_ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__and2_1
XFILLER_38_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13480_ _06162_ _06236_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__nand2_1
X_10692_ _03483_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__buf_6
XFILLER_185_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12431_ _05133_ _05147_ _05187_ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__o21ai_2
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15150_ _07265_ _07332_ _07786_ _06873_ vssd1 vssd1 vccd1 vccd1 _07837_ sky130_fd_sc_hd__o22ai_1
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12362_ _05116_ _05118_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__or2_1
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14101_ rbzero.wall_tracer.trackDistX\[10\] rbzero.wall_tracer.trackDistY\[10\] _06783_
+ vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__a21o_1
XFILLER_153_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11313_ rbzero.debug_overlay.vplaneX\[-7\] _04083_ _04084_ rbzero.debug_overlay.vplaneX\[-6\]
+ gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__a221o_1
X_15081_ _07765_ _07767_ _07187_ _07768_ vssd1 vssd1 vccd1 vccd1 _07769_ sky130_fd_sc_hd__o31a_1
X_12293_ _05049_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__inv_2
XFILLER_10_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14032_ _06769_ _06770_ _06630_ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__a21oi_4
X_11244_ _03860_ _04018_ _04028_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__and3b_1
XFILLER_101_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11175_ rbzero.tex_r1\[7\] _03925_ _03959_ _03726_ vssd1 vssd1 vccd1 vccd1 _03960_
+ sky130_fd_sc_hd__o211a_1
X_18840_ rbzero.pov.ready_buffer\[1\] _02663_ _02682_ _02672_ vssd1 vssd1 vccd1 vccd1
+ _01060_ sky130_fd_sc_hd__o211a_1
XFILLER_171_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10126_ rbzero.tex_g1\[4\] rbzero.tex_g1\[5\] _03117_ vssd1 vssd1 vccd1 vccd1 _03121_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__02440_ _02440_ vssd1 vssd1 vccd1 vccd1 clknet_0__02440_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18771_ _02638_ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15983_ _08199_ _08314_ vssd1 vssd1 vccd1 vccd1 _08597_ sky130_fd_sc_hd__nor2_1
XFILLER_121_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17722_ rbzero.debug_overlay.vplaneX\[-3\] rbzero.debug_overlay.vplaneX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__and2_1
X_14934_ _07589_ _07592_ vssd1 vssd1 vccd1 vccd1 _07622_ sky130_fd_sc_hd__xnor2_1
X_10057_ rbzero.tex_g1\[37\] rbzero.tex_g1\[38\] _03084_ vssd1 vssd1 vccd1 vccd1 _03085_
+ sky130_fd_sc_hd__mux2_1
XFILLER_169_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17653_ _01918_ _01929_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14865_ _07504_ _07507_ vssd1 vssd1 vccd1 vccd1 _07553_ sky130_fd_sc_hd__xnor2_2
XFILLER_180_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16604_ _09150_ _09212_ vssd1 vssd1 vccd1 vccd1 _09213_ sky130_fd_sc_hd__nand2_2
XFILLER_169_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13816_ _06569_ _06284_ vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__and2b_1
X_17584_ _01863_ _01864_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__or2_1
XFILLER_51_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14796_ _06893_ _06917_ _06954_ _06977_ vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__or4_1
X_19226__382 clknet_1_1__leaf__02753_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__inv_2
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19323_ rbzero.texV\[-1\] _02762_ _02709_ _02809_ vssd1 vssd1 vccd1 vccd1 _01416_
+ sky130_fd_sc_hd__a22o_1
X_16535_ _09021_ _09133_ _09018_ _09015_ vssd1 vssd1 vccd1 vccd1 _09145_ sky130_fd_sc_hd__o31a_1
XFILLER_16_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13747_ _06496_ _06502_ _06503_ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__nand3b_1
X_10959_ _03674_ _03738_ _03744_ _03704_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__a211o_1
XFILLER_31_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16466_ _08952_ _08953_ vssd1 vssd1 vccd1 vccd1 _09077_ sky130_fd_sc_hd__nand2_1
XFILLER_32_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13678_ _06382_ _06425_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__xnor2_2
X_18205_ rbzero.color_sky\[1\] rbzero.spi_registers.new_sky\[1\] _02320_ vssd1 vssd1
+ vccd1 vccd1 _02324_ sky130_fd_sc_hd__mux2_1
X_15417_ _07039_ _07141_ vssd1 vssd1 vccd1 vccd1 _08102_ sky130_fd_sc_hd__or2_1
X_12629_ _05215_ _05305_ _05302_ _05306_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__or4_1
X_16397_ _09007_ _08896_ vssd1 vssd1 vccd1 vccd1 _09008_ sky130_fd_sc_hd__nor2_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18136_ _03467_ _03503_ _03911_ _03505_ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__and4b_1
XFILLER_156_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15348_ _07886_ _07909_ _08033_ vssd1 vssd1 vccd1 vccd1 _08034_ sky130_fd_sc_hd__a21oi_1
XFILLER_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18067_ _02237_ vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15279_ _07871_ _07942_ _07963_ vssd1 vssd1 vccd1 vccd1 _07965_ sky130_fd_sc_hd__nand3_1
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17018_ rbzero.wall_tracer.trackDistX\[8\] rbzero.wall_tracer.stepDistX\[8\] vssd1
+ vssd1 vccd1 vccd1 _09624_ sky130_fd_sc_hd__nand2_1
XFILLER_172_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09840_ rbzero.tex_r1\[10\] rbzero.tex_r1\[11\] _02965_ vssd1 vssd1 vccd1 vccd1 _02969_
+ sky130_fd_sc_hd__mux2_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ rbzero.tex_r1\[43\] rbzero.tex_r1\[44\] _02932_ vssd1 vssd1 vccd1 vccd1 _02933_
+ sky130_fd_sc_hd__mux2_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20227_ net287 _01158_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[10\] sky130_fd_sc_hd__dfxtp_1
X_20158_ net218 _01089_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09969_ rbzero.tex_r0\[15\] rbzero.tex_r0\[14\] _03028_ vssd1 vssd1 vccd1 vccd1 _03038_
+ sky130_fd_sc_hd__mux2_1
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12980_ _05526_ _05433_ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__nor2_1
X_20089_ clknet_leaf_8_i_clk _01020_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11931_ _04672_ _03913_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__nor2_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _07336_ _07337_ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__nor2_2
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _04631_ _04636_ _04637_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__o21ai_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _06309_ _06321_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__xnor2_1
X_10813_ _03583_ _03598_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__nor2_1
XFILLER_14_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _06873_ vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__buf_2
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18394__37 clknet_1_0__leaf__02435_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__inv_2
X_11793_ net16 net15 vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__and2_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16320_ _08922_ _08931_ vssd1 vssd1 vccd1 vccd1 _08932_ sky130_fd_sc_hd__xnor2_1
X_13532_ _06288_ vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10744_ _03461_ _03467_ _03525_ _03529_ _02902_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__o41a_1
XFILLER_201_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16251_ _07012_ _08862_ _08359_ vssd1 vssd1 vccd1 vccd1 _08863_ sky130_fd_sc_hd__or3_1
XFILLER_201_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13463_ _06202_ _06203_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__nor2_1
XFILLER_90_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10675_ _02902_ _03468_ _03469_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__o21ai_1
XFILLER_90_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15202_ _07661_ _07766_ _07748_ _07662_ vssd1 vssd1 vccd1 vccd1 _07889_ sky130_fd_sc_hd__o22ai_1
XFILLER_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12414_ _05062_ _05060_ _05061_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__a21o_1
X_16182_ _08788_ _08793_ vssd1 vssd1 vccd1 vccd1 _08795_ sky130_fd_sc_hd__or2_1
XFILLER_127_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13394_ _06149_ _06150_ vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15133_ _07813_ _07814_ _07820_ vssd1 vssd1 vccd1 vccd1 _07821_ sky130_fd_sc_hd__a21oi_1
X_12345_ _05100_ _05101_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__xnor2_2
XFILLER_182_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19941_ net170 _00872_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[21\] sky130_fd_sc_hd__dfxtp_1
X_15064_ _04831_ _07750_ _07751_ _07162_ vssd1 vssd1 vccd1 vccd1 _07752_ sky130_fd_sc_hd__a31o_1
X_12276_ rbzero.debug_overlay.facingX\[-4\] rbzero.wall_tracer.rayAddendX\[4\] vssd1
+ vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__nor2_1
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14015_ _05334_ _06703_ _06755_ _06756_ _05369_ vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__o221a_1
X_11227_ _03834_ _03517_ _03908_ _04011_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__a31o_1
XFILLER_96_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19872_ clknet_leaf_21_i_clk _00803_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18823_ rbzero.pov.ready_buffer\[15\] _02666_ _02673_ _02651_ vssd1 vssd1 vccd1 vccd1
+ _01052_ sky130_fd_sc_hd__a211o_1
XFILLER_68_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11158_ rbzero.tex_r1\[44\] _03920_ _03925_ _03941_ _03942_ vssd1 vssd1 vccd1 vccd1
+ _03943_ sky130_fd_sc_hd__a311o_1
XFILLER_95_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10109_ rbzero.tex_g1\[12\] rbzero.tex_g1\[13\] _03106_ vssd1 vssd1 vccd1 vccd1 _03112_
+ sky130_fd_sc_hd__mux2_1
XFILLER_191_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18754_ _02628_ _02631_ _02559_ vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__a21oi_1
X_11089_ _03840_ rbzero.map_overlay.i_othery\[4\] rbzero.map_overlay.i_otherx\[2\]
+ _03781_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__a22o_1
X_15966_ _08578_ _08579_ _08580_ vssd1 vssd1 vccd1 vccd1 _08582_ sky130_fd_sc_hd__a21o_1
XFILLER_110_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14917_ _07584_ _07604_ vssd1 vssd1 vccd1 vccd1 _07605_ sky130_fd_sc_hd__or2_1
X_17705_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.debug_overlay.vplaneX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__or2_1
X_18685_ _02543_ _02576_ rbzero.debug_overlay.playerX\[5\] vssd1 vssd1 vccd1 vccd1
+ _02578_ sky130_fd_sc_hd__a21boi_1
X_15897_ _08518_ _08519_ _08513_ vssd1 vssd1 vccd1 vccd1 _08521_ sky130_fd_sc_hd__a21bo_1
X_14848_ _07531_ _07535_ _07534_ vssd1 vssd1 vccd1 vccd1 _07536_ sky130_fd_sc_hd__a21oi_1
XFILLER_24_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17636_ rbzero.debug_overlay.playerY\[5\] _01913_ _09620_ vssd1 vssd1 vccd1 vccd1
+ _01914_ sky130_fd_sc_hd__mux2_1
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17567_ _01785_ rbzero.wall_tracer.rayAddendY\[7\] vssd1 vssd1 vccd1 vccd1 _01854_
+ sky130_fd_sc_hd__or2_1
X_14779_ _07463_ _07465_ _07466_ vssd1 vssd1 vccd1 vccd1 _07467_ sky130_fd_sc_hd__a21oi_1
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16518_ _09027_ _09099_ _09126_ vssd1 vssd1 vccd1 vccd1 _09128_ sky130_fd_sc_hd__nand3_1
X_19306_ rbzero.traced_texa\[-3\] rbzero.texV\[-3\] vssd1 vssd1 vccd1 vccd1 _02795_
+ sky130_fd_sc_hd__and2_1
XFILLER_147_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17498_ _04109_ rbzero.debug_overlay.vplaneY\[-6\] vssd1 vssd1 vccd1 vccd1 _01790_
+ sky130_fd_sc_hd__xor2_1
XFILLER_56_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16449_ _09058_ _09059_ vssd1 vssd1 vccd1 vccd1 _09060_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18119_ rbzero.spi_registers.new_other\[8\] _02264_ _02269_ _02266_ vssd1 vssd1 vccd1
+ vccd1 _00752_ sky130_fd_sc_hd__o211a_1
XFILLER_172_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20012_ clknet_leaf_91_i_clk _00943_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09823_ rbzero.tex_r1\[18\] rbzero.tex_r1\[19\] _02954_ vssd1 vssd1 vccd1 vccd1 _02960_
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09754_ rbzero.tex_r1\[51\] rbzero.tex_r1\[52\] _02921_ vssd1 vssd1 vccd1 vccd1 _02924_
+ sky130_fd_sc_hd__mux2_1
XFILLER_101_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10460_ rbzero.tex_b0\[38\] rbzero.tex_b0\[37\] _03291_ vssd1 vssd1 vccd1 vccd1 _03296_
+ sky130_fd_sc_hd__mux2_1
XFILLER_195_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10391_ rbzero.tex_b1\[6\] rbzero.tex_b1\[7\] _03254_ vssd1 vssd1 vccd1 vccd1 _03260_
+ sky130_fd_sc_hd__mux2_1
XFILLER_191_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18919__105 clknet_1_0__leaf__02723_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__inv_2
XFILLER_191_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12130_ _04857_ _04891_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__nand2_1
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12061_ _04830_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__clkbuf_4
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11012_ rbzero.row_render.size\[7\] _03775_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15820_ _08458_ vssd1 vssd1 vccd1 vccd1 _08462_ sky130_fd_sc_hd__clkbuf_4
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _08431_ _08433_ vssd1 vssd1 vccd1 vccd1 _08434_ sky130_fd_sc_hd__xnor2_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12963_ _05700_ _05719_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__nor2_1
XFILLER_92_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _07383_ _07389_ vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__xnor2_1
XFILLER_166_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18470_ _02451_ vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11914_ clknet_1_0__leaf__04486_ _04668_ _04685_ _04686_ _04688_ vssd1 vssd1 vccd1
+ vccd1 _04689_ sky130_fd_sc_hd__a311o_2
XFILLER_166_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15682_ _08229_ _07878_ vssd1 vssd1 vccd1 vccd1 _08365_ sky130_fd_sc_hd__nor2_1
XFILLER_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _05494_ _05576_ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__nand2_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _01716_ _01717_ _01718_ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__or3_1
XFILLER_33_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _07259_ _07260_ vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__or2_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ net12 _04614_ _04618_ _04620_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__o211a_1
XFILLER_54_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _01668_ vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14564_ _07042_ _07049_ _07052_ _07041_ vssd1 vssd1 vccd1 vccd1 _07252_ sky130_fd_sc_hd__o31a_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _04552_ _03913_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__nor2_1
XFILLER_159_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16303_ _06997_ _08134_ vssd1 vssd1 vccd1 vccd1 _08915_ sky130_fd_sc_hd__nor2_1
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13515_ _06253_ _06270_ _06271_ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__a21oi_1
X_10727_ gpout0.hpos\[7\] _03512_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__and2_1
X_17283_ _01609_ _01610_ _01611_ vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__and3_1
XFILLER_201_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14495_ rbzero.wall_tracer.visualWallDist\[-10\] _04841_ _06860_ _07152_ vssd1 vssd1
+ vccd1 vccd1 _07183_ sky130_fd_sc_hd__and4_1
XFILLER_146_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16234_ _08844_ _08845_ vssd1 vssd1 vccd1 vccd1 _08846_ sky130_fd_sc_hd__nor2_1
XFILLER_146_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13446_ _06102_ _06112_ _06114_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__o21a_1
X_10658_ _03404_ _03450_ _03453_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__and3_1
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16165_ _08108_ _07878_ _08649_ _08648_ vssd1 vssd1 vccd1 vccd1 _08778_ sky130_fd_sc_hd__o31a_1
XFILLER_127_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13377_ _06120_ _06133_ _06132_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__a21oi_1
X_19037__211 clknet_1_1__leaf__02735_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__inv_2
X_10589_ rbzero.wall_tracer.visualWallDist\[3\] rbzero.wall_tracer.visualWallDist\[2\]
+ rbzero.wall_tracer.visualWallDist\[1\] rbzero.wall_tracer.visualWallDist\[0\] vssd1
+ vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__or4_1
XFILLER_115_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15116_ _07076_ _07371_ _07369_ vssd1 vssd1 vccd1 vccd1 _07804_ sky130_fd_sc_hd__a21o_2
X_12328_ _05052_ _05083_ _05084_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__a21bo_1
XFILLER_141_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16096_ _08598_ _08709_ vssd1 vssd1 vccd1 vccd1 _08710_ sky130_fd_sc_hd__xor2_1
XFILLER_6_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15047_ _07078_ vssd1 vssd1 vccd1 vccd1 _07735_ sky130_fd_sc_hd__buf_2
X_19924_ net153 _00855_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[4\] sky130_fd_sc_hd__dfxtp_1
X_12259_ _05017_ _05018_ rbzero.wall_tracer.mapY\[8\] _05009_ vssd1 vssd1 vccd1 vccd1
+ _00403_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_123_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19855_ clknet_leaf_21_i_clk _00786_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_18806_ rbzero.debug_overlay.facingY\[-1\] _02660_ vssd1 vssd1 vccd1 vccd1 _02664_
+ sky130_fd_sc_hd__or2_1
XFILLER_95_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19786_ clknet_leaf_86_i_clk _00717_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[68\]
+ sky130_fd_sc_hd__dfxtp_1
X_16998_ _09531_ _09603_ vssd1 vssd1 vccd1 vccd1 _09604_ sky130_fd_sc_hd__nand2_1
XFILLER_77_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18737_ rbzero.debug_overlay.playerY\[2\] _02588_ _02617_ _02586_ vssd1 vssd1 vccd1
+ vccd1 _01022_ sky130_fd_sc_hd__o211a_1
XFILLER_95_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15949_ _08563_ _08564_ _08565_ vssd1 vssd1 vccd1 vccd1 _08567_ sky130_fd_sc_hd__a21o_1
XFILLER_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18668_ rbzero.pov.ready_buffer\[69\] _02411_ _02535_ _02564_ _02543_ vssd1 vssd1
+ vccd1 vccd1 _02565_ sky130_fd_sc_hd__o221a_1
X_19083__253 clknet_1_0__leaf__02739_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__inv_2
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17619_ _04936_ _04939_ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__xor2_1
XFILLER_52_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18599_ rbzero.pov.spi_buffer\[67\] rbzero.pov.spi_buffer\[68\] _02510_ vssd1 vssd1
+ vccd1 vccd1 _02519_ sky130_fd_sc_hd__mux2_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20492_ clknet_leaf_43_i_clk _01423_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09806_ rbzero.tex_r1\[26\] rbzero.tex_r1\[27\] _02943_ vssd1 vssd1 vccd1 vccd1 _02951_
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09737_ rbzero.tex_r1\[59\] rbzero.tex_r1\[60\] _02910_ vssd1 vssd1 vccd1 vccd1 _02915_
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18451__88 clknet_1_0__leaf__02441_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__inv_2
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ rbzero.tex_b1\[33\] rbzero.tex_b1\[32\] _03616_ vssd1 vssd1 vccd1 vccd1 _04411_
+ sky130_fd_sc_hd__mux2_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11561_ rbzero.tex_b0\[41\] rbzero.tex_b0\[40\] _04188_ vssd1 vssd1 vccd1 vccd1 _04343_
+ sky130_fd_sc_hd__mux2_1
XFILLER_129_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13300_ _05549_ _05576_ _06056_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__and3_1
X_10512_ rbzero.tex_b0\[13\] rbzero.tex_b0\[12\] _03313_ vssd1 vssd1 vccd1 vccd1 _03323_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14280_ _06949_ vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__clkbuf_4
X_11492_ rbzero.tex_g1\[49\] rbzero.tex_g1\[48\] _04247_ vssd1 vssd1 vccd1 vccd1 _04275_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13231_ _05987_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__clkbuf_4
XFILLER_108_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10443_ rbzero.tex_b0\[46\] rbzero.tex_b0\[45\] _03280_ vssd1 vssd1 vccd1 vccd1 _03287_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18911__97 clknet_1_1__leaf__02723_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__inv_2
XFILLER_152_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13162_ _05469_ _05918_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__xor2_1
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10374_ rbzero.tex_b1\[14\] rbzero.tex_b1\[15\] _03243_ vssd1 vssd1 vccd1 vccd1 _03251_
+ sky130_fd_sc_hd__mux2_1
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12113_ _04870_ _04874_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__or2b_1
XFILLER_112_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17970_ _02185_ vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__clkbuf_1
X_13093_ _05760_ _05800_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__and2b_1
X_16921_ _09372_ _09431_ _09459_ vssd1 vssd1 vccd1 vccd1 _09527_ sky130_fd_sc_hd__a21o_1
XFILLER_137_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12044_ _04787_ _04816_ net34 net35 vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__o211a_1
XFILLER_77_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19640_ clknet_leaf_39_i_clk _00571_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16852_ _09443_ _09458_ vssd1 vssd1 vccd1 vccd1 _09459_ sky130_fd_sc_hd__xnor2_1
XFILLER_78_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15803_ rbzero.row_render.texu\[5\] _08457_ _08453_ rbzero.wall_tracer.texu\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__a22o_1
X_16783_ _09375_ _09390_ vssd1 vssd1 vccd1 vccd1 _09391_ sky130_fd_sc_hd__nand2_1
X_19571_ clknet_leaf_36_i_clk _00502_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13995_ _06739_ vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__clkbuf_1
X_15734_ _08356_ _08284_ _08416_ vssd1 vssd1 vccd1 vccd1 _08417_ sky130_fd_sc_hd__a21oi_1
X_18522_ rbzero.pov.spi_buffer\[30\] rbzero.pov.spi_buffer\[31\] _02477_ vssd1 vssd1
+ vccd1 vccd1 _02479_ sky130_fd_sc_hd__mux2_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12946_ _05667_ _05702_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15665_ _08346_ _08347_ vssd1 vssd1 vccd1 vccd1 _08348_ sky130_fd_sc_hd__nor2_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ _05473_ _05517_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__or2_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ rbzero.debug_overlay.vplaneY\[-6\] rbzero.wall_tracer.rayAddendY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__or2_1
XFILLER_61_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _06900_ _06933_ vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__nor2_1
X_11828_ _03852_ _04552_ net17 _04604_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__a211o_1
X_15596_ _08278_ _08279_ vssd1 vssd1 vccd1 vccd1 _08280_ sky130_fd_sc_hd__nor2_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _08485_ _01655_ _01656_ _01522_ vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__o31a_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _06969_ vssd1 vssd1 vccd1 vccd1 _07235_ sky130_fd_sc_hd__clkbuf_4
XFILLER_105_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11759_ _04522_ _04535_ _04514_ net42 _04536_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__a221o_1
XFILLER_147_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17266_ rbzero.wall_tracer.trackDistY\[0\] rbzero.wall_tracer.stepDistY\[0\] _01592_
+ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__a21o_1
X_14478_ _07163_ _07164_ _07165_ _04831_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__o211a_1
X_16217_ _08601_ _08828_ vssd1 vssd1 vccd1 vccd1 _08830_ sky130_fd_sc_hd__or2_1
XFILLER_174_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13429_ _06183_ _06185_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__nand2_1
XFILLER_174_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17197_ _01535_ _01536_ _01537_ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__or3_1
XFILLER_127_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16148_ _08657_ _08729_ _08759_ vssd1 vssd1 vccd1 vccd1 _08761_ sky130_fd_sc_hd__nand3_1
XFILLER_170_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16079_ _08671_ _08692_ vssd1 vssd1 vccd1 vccd1 _08693_ sky130_fd_sc_hd__xnor2_2
X_19907_ clknet_leaf_24_i_clk _00838_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19838_ clknet_leaf_15_i_clk _00769_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_110_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 i_debug_map_overlay vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_4
X_19769_ clknet_leaf_6_i_clk _00700_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_18948__131 clknet_1_1__leaf__02726_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__inv_2
XFILLER_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20475_ clknet_leaf_37_i_clk _01406_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18994__173 clknet_1_0__leaf__02730_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__inv_2
XFILLER_195_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10090_ rbzero.tex_g1\[21\] rbzero.tex_g1\[22\] _03095_ vssd1 vssd1 vccd1 vccd1 _03102_
+ sky130_fd_sc_hd__mux2_1
XFILLER_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_7_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12800_ _05416_ _05417_ _05424_ _05210_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__and4b_2
XFILLER_28_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13780_ _06383_ _06536_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__nand2_1
X_10992_ rbzero.row_render.size\[7\] rbzero.row_render.size\[6\] rbzero.row_render.size\[8\]
+ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__a21o_1
XFILLER_43_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12731_ _05443_ _05404_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__nor2_4
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15450_ _07661_ _08133_ _08134_ _07662_ vssd1 vssd1 vccd1 vccd1 _08135_ sky130_fd_sc_hd__o22ai_1
XFILLER_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _05383_ _05386_ _05338_ vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__a21o_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _04830_ _07088_ vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__or2_1
XFILLER_187_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11613_ rbzero.color_sky\[5\] rbzero.color_floor\[5\] _03535_ vssd1 vssd1 vccd1 vccd1
+ _04394_ sky130_fd_sc_hd__mux2_1
X_15381_ _07958_ _07962_ _07956_ vssd1 vssd1 vccd1 vccd1 _08066_ sky130_fd_sc_hd__a21o_1
XFILLER_11_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12593_ _05178_ _05223_ _05349_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__mux2_1
XFILLER_184_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17120_ _08862_ _08317_ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__nand2_1
X_14332_ rbzero.wall_tracer.visualWallDist\[-2\] _06985_ _06906_ vssd1 vssd1 vccd1
+ vccd1 _07020_ sky130_fd_sc_hd__a21oi_1
XFILLER_196_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11544_ _04324_ _04325_ _03660_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__mux2_1
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17051_ _09633_ _09654_ _09655_ _09653_ vssd1 vssd1 vccd1 vccd1 _09656_ sky130_fd_sc_hd__o22a_1
XFILLER_51_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14263_ rbzero.wall_tracer.side _04894_ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__nor2_1
XFILLER_52_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11475_ rbzero.tex_g1\[14\] _03618_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__and2_1
XFILLER_143_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16002_ _08339_ vssd1 vssd1 vccd1 vccd1 _08616_ sky130_fd_sc_hd__inv_2
XFILLER_183_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__02740_ _02740_ vssd1 vssd1 vccd1 vccd1 clknet_0__02740_ sky130_fd_sc_hd__clkbuf_16
X_13214_ _05959_ _05970_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__xnor2_1
XFILLER_109_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10426_ rbzero.tex_b0\[54\] rbzero.tex_b0\[53\] _03269_ vssd1 vssd1 vccd1 vccd1 _03278_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14194_ rbzero.wall_tracer.rayAddendX\[-3\] rbzero.wall_tracer.rayAddendX\[-2\] _05113_
+ _05107_ vssd1 vssd1 vccd1 vccd1 _06882_ sky130_fd_sc_hd__or4_1
XFILLER_136_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13145_ _05836_ _05847_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__xnor2_2
X_10357_ rbzero.tex_b1\[22\] rbzero.tex_b1\[23\] _03232_ vssd1 vssd1 vccd1 vccd1 _03242_
+ sky130_fd_sc_hd__mux2_1
XFILLER_140_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _05796_ _05791_ _05795_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__or3_1
X_17953_ rbzero.pov.spi_buffer\[30\] rbzero.pov.ready_buffer\[30\] _02175_ vssd1 vssd1
+ vccd1 vccd1 _02177_ sky130_fd_sc_hd__mux2_1
X_10288_ rbzero.tex_b1\[55\] rbzero.tex_b1\[56\] _03199_ vssd1 vssd1 vccd1 vccd1 _03206_
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16904_ _09508_ _09510_ vssd1 vssd1 vccd1 vccd1 _09511_ sky130_fd_sc_hd__nor2_1
X_12027_ net49 net40 net39 _03537_ net34 _04790_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__mux4_1
XFILLER_78_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19149__312 clknet_1_1__leaf__02746_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__inv_2
X_17884_ _02139_ vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19623_ clknet_leaf_48_i_clk _00554_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16835_ _09439_ _09440_ vssd1 vssd1 vccd1 vccd1 _09442_ sky130_fd_sc_hd__or2_1
XFILLER_65_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19554_ clknet_leaf_9_i_clk _00485_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[4\] sky130_fd_sc_hd__dfxtp_2
X_16766_ _09372_ _09373_ vssd1 vssd1 vccd1 vccd1 _09374_ sky130_fd_sc_hd__nand2_1
X_13978_ _05390_ _06724_ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__nor2_1
XFILLER_93_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18505_ rbzero.pov.spi_buffer\[22\] rbzero.pov.spi_buffer\[23\] _02466_ vssd1 vssd1
+ vccd1 vccd1 _02470_ sky130_fd_sc_hd__mux2_1
X_15717_ _03388_ _07185_ _08396_ _08399_ vssd1 vssd1 vccd1 vccd1 _08400_ sky130_fd_sc_hd__or4_1
X_12929_ _05664_ _05684_ _05685_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__a21boi_1
X_16697_ _09305_ _09196_ vssd1 vssd1 vccd1 vccd1 _09306_ sky130_fd_sc_hd__and2_1
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19485_ clknet_leaf_57_i_clk _00431_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_61_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15648_ _08328_ _08329_ vssd1 vssd1 vccd1 vccd1 _08331_ sky130_fd_sc_hd__nand2_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15579_ _07877_ _08133_ vssd1 vssd1 vccd1 vccd1 _08263_ sky130_fd_sc_hd__nor2_1
X_18367_ rbzero.pov.spi_counter\[2\] _02417_ _02415_ vssd1 vssd1 vccd1 vccd1 _02424_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_159_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17318_ _01634_ _01637_ _01635_ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__o21ai_1
XFILLER_186_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19195__354 clknet_1_0__leaf__02750_ vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__inv_2
X_18298_ _02382_ vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17249_ _01534_ _01581_ _01582_ _01526_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__a31o_1
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20260_ net320 _01191_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20191_ net251 _01122_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19015__191 clknet_1_1__leaf__02733_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__inv_2
XFILLER_116_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_50 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_61 _08958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_72 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11260_ _04037_ _04044_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__or2_1
XFILLER_197_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20458_ net138 _01389_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10211_ _03165_ vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11191_ _03648_ _03971_ _03975_ _03687_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__a31o_1
X_20389_ net449 _01320_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10142_ rbzero.tex_g0\[61\] rbzero.tex_g0\[60\] _03050_ vssd1 vssd1 vccd1 vccd1 _03129_
+ sky130_fd_sc_hd__mux2_1
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14950_ _07541_ _07632_ _07637_ vssd1 vssd1 vccd1 vccd1 _07638_ sky130_fd_sc_hd__or3_1
X_10073_ rbzero.tex_g1\[29\] rbzero.tex_g1\[30\] _03084_ vssd1 vssd1 vccd1 vccd1 _03093_
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13901_ _05421_ _06655_ _06613_ _05372_ _06637_ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__o221a_1
XFILLER_130_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14881_ _07545_ _07567_ vssd1 vssd1 vccd1 vccd1 _07569_ sky130_fd_sc_hd__or2b_1
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16620_ _07787_ vssd1 vssd1 vccd1 vccd1 _09229_ sky130_fd_sc_hd__buf_2
X_13832_ _06572_ _06587_ _06588_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__mux2_1
XFILLER_90_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16551_ _09048_ _09155_ _09160_ vssd1 vssd1 vccd1 vccd1 _09161_ sky130_fd_sc_hd__a21o_1
XFILLER_16_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13763_ _06487_ _06519_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__xor2_1
X_10975_ _03666_ _03758_ _03759_ _03760_ _03702_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__o221a_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15502_ _08092_ _08066_ vssd1 vssd1 vccd1 vccd1 _08186_ sky130_fd_sc_hd__or2b_1
X_12714_ _05470_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__buf_2
X_16482_ _09078_ _09089_ _09090_ _08957_ _09091_ vssd1 vssd1 vccd1 vccd1 _09092_ sky130_fd_sc_hd__a221o_1
X_19270_ _02763_ _02764_ _02760_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__a21bo_1
X_13694_ _06406_ _06415_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__xor2_1
XFILLER_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15433_ _07581_ _07198_ vssd1 vssd1 vccd1 vccd1 _08118_ sky130_fd_sc_hd__nor2_1
XFILLER_31_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18221_ rbzero.spi_registers.got_new_floor _02261_ vssd1 vssd1 vccd1 vccd1 _02335_
+ sky130_fd_sc_hd__and2_2
X_12645_ _05330_ _05377_ _05371_ _05325_ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_54_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15364_ _07703_ _07807_ _07927_ vssd1 vssd1 vccd1 vccd1 _08050_ sky130_fd_sc_hd__a21oi_1
XFILLER_15_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18152_ rbzero.spi_registers.new_mapd\[10\] _02290_ _02293_ _02275_ vssd1 vssd1 vccd1
+ vccd1 _00761_ sky130_fd_sc_hd__o211a_1
X_12576_ _05321_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__clkbuf_4
XFILLER_156_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17103_ _09706_ _09707_ _08509_ vssd1 vssd1 vccd1 vccd1 _09708_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14315_ _06850_ _05107_ _07002_ _04830_ vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__a211o_1
XFILLER_184_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18083_ _02246_ vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__clkbuf_1
X_11527_ _04028_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__inv_2
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15295_ _07860_ _07979_ _07980_ vssd1 vssd1 vccd1 vccd1 _07981_ sky130_fd_sc_hd__o21bai_1
XFILLER_144_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17034_ _09541_ _09637_ _09638_ vssd1 vssd1 vccd1 vccd1 _09639_ sky130_fd_sc_hd__a21bo_1
XFILLER_171_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14246_ _03490_ rbzero.wall_tracer.stepDistY\[-5\] rbzero.wall_tracer.state\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__a21o_1
XFILLER_109_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11458_ rbzero.tex_g1\[17\] rbzero.tex_g1\[16\] _03700_ vssd1 vssd1 vccd1 vccd1 _04241_
+ sky130_fd_sc_hd__mux2_1
XFILLER_144_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__02723_ _02723_ vssd1 vssd1 vccd1 vccd1 clknet_0__02723_ sky130_fd_sc_hd__clkbuf_16
X_10409_ _03143_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__clkbuf_4
X_14177_ _04949_ rbzero.wall_tracer.stepDistX\[-11\] _06864_ vssd1 vssd1 vccd1 vccd1
+ _06865_ sky130_fd_sc_hd__a21oi_4
X_11389_ rbzero.tex_g0\[3\] rbzero.tex_g0\[2\] _03615_ vssd1 vssd1 vccd1 vccd1 _04173_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13128_ _05877_ _05884_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__xnor2_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17936_ rbzero.pov.spi_buffer\[22\] rbzero.pov.ready_buffer\[22\] _02164_ vssd1 vssd1
+ vccd1 vccd1 _02168_ sky130_fd_sc_hd__mux2_1
X_13059_ _05809_ _05815_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__and2_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17867_ rbzero.spi_registers.spi_counter\[2\] _02112_ _02122_ vssd1 vssd1 vccd1 vccd1
+ _02126_ sky130_fd_sc_hd__o21ai_1
X_19606_ clknet_leaf_63_i_clk _00537_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_16818_ _09332_ _09333_ _09330_ vssd1 vssd1 vccd1 vccd1 _09425_ sky130_fd_sc_hd__a21oi_1
XFILLER_94_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17798_ _02000_ rbzero.wall_tracer.rayAddendX\[7\] vssd1 vssd1 vccd1 vccd1 _02063_
+ sky130_fd_sc_hd__or2_1
XFILLER_35_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19537_ clknet_leaf_62_i_clk _00008_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_16749_ _09009_ _09007_ _09142_ _08134_ vssd1 vssd1 vccd1 vccd1 _09357_ sky130_fd_sc_hd__or4_1
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19468_ clknet_leaf_61_i_clk _00414_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19203__361 clknet_1_0__leaf__02751_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__inv_2
XFILLER_166_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19399_ rbzero.traced_texVinit\[5\] _02868_ _08174_ _01745_ vssd1 vssd1 vccd1 vccd1
+ _01433_ sky130_fd_sc_hd__a22o_1
XFILLER_107_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20312_ net372 _01243_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20243_ net303 _01174_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20174_ net234 _01105_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09985_ _03046_ vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_72_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_87_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_199_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10760_ _03544_ _03545_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__nand2_1
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_10691_ rbzero.vga_sync.vsync _02981_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__nor2_2
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12430_ _03489_ _05078_ _05151_ _05080_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__o31ai_2
XFILLER_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12361_ rbzero.wall_tracer.rayAddendX\[-2\] _05117_ _05072_ vssd1 vssd1 vccd1 vccd1
+ _05118_ sky130_fd_sc_hd__mux2_2
XFILLER_193_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14100_ rbzero.wall_tracer.visualWallDist\[9\] _03496_ _06814_ _03498_ vssd1 vssd1
+ vccd1 vccd1 _00448_ sky130_fd_sc_hd__o211a_1
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11312_ rbzero.debug_overlay.facingY\[-2\] _04056_ _04096_ vssd1 vssd1 vccd1 vccd1
+ _04097_ sky130_fd_sc_hd__a21oi_1
X_15080_ _07143_ _07188_ vssd1 vssd1 vccd1 vccd1 _07768_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_25_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12292_ _05031_ _05035_ _05033_ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__a21o_1
XFILLER_154_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14031_ _05315_ _06750_ _06763_ _05373_ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__a31o_1
X_11243_ _03838_ _04019_ _04022_ _04027_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__a31o_1
XFILLER_180_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11174_ rbzero.tex_r1\[6\] _03926_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__or2_1
X_19031__206 clknet_1_0__leaf__02734_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__inv_2
XFILLER_161_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10125_ _03120_ vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18770_ rbzero.pov.ready_buffer\[36\] _02636_ _02642_ _02643_ vssd1 vssd1 vccd1 vccd1
+ _01029_ sky130_fd_sc_hd__o211a_1
X_15982_ _08594_ _08589_ _08592_ _08593_ vssd1 vssd1 vccd1 vccd1 _08596_ sky130_fd_sc_hd__a211oi_2
X_17721_ rbzero.debug_overlay.vplaneX\[-3\] rbzero.debug_overlay.vplaneX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__nor2_1
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14933_ _07616_ _07620_ vssd1 vssd1 vccd1 vccd1 _07621_ sky130_fd_sc_hd__xnor2_1
X_10056_ _03072_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__clkbuf_4
X_17652_ _01919_ _01927_ _01928_ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__a21boi_1
XFILLER_169_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14864_ _07531_ _07535_ vssd1 vssd1 vccd1 vccd1 _07552_ sky130_fd_sc_hd__xor2_1
XFILLER_29_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16603_ _09152_ _09131_ vssd1 vssd1 vccd1 vccd1 _09212_ sky130_fd_sc_hd__or2b_1
X_13815_ _06211_ _06571_ vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__xor2_2
X_14795_ _07119_ _06978_ vssd1 vssd1 vccd1 vccd1 _07483_ sky130_fd_sc_hd__nor2_1
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17583_ _01853_ _01858_ _01867_ _03339_ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__a31o_1
XFILLER_189_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19322_ _02807_ _02808_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__xor2_1
X_16534_ _09141_ _09143_ vssd1 vssd1 vccd1 vccd1 _09144_ sky130_fd_sc_hd__xor2_1
X_13746_ _06461_ _06479_ _06495_ vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__a21o_1
XFILLER_189_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10958_ _03740_ _03741_ _03743_ _03670_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__o211a_1
XFILLER_91_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16465_ _08967_ _09075_ vssd1 vssd1 vccd1 vccd1 _09076_ sky130_fd_sc_hd__xor2_2
XFILLER_32_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13677_ _06335_ _06433_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__xnor2_1
X_10889_ rbzero.tex_r0\[9\] rbzero.tex_r0\[8\] _03663_ vssd1 vssd1 vccd1 vccd1 _03675_
+ sky130_fd_sc_hd__mux2_1
XFILLER_189_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18204_ _04827_ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__clkbuf_4
X_15416_ _08099_ _08100_ vssd1 vssd1 vccd1 vccd1 _08101_ sky130_fd_sc_hd__xnor2_1
X_12628_ _05383_ _05384_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__nand2_1
X_16396_ _07012_ vssd1 vssd1 vccd1 vccd1 _09007_ sky130_fd_sc_hd__buf_2
XFILLER_192_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15347_ _07906_ _07908_ vssd1 vssd1 vccd1 vccd1 _08033_ sky130_fd_sc_hd__nor2_1
X_18135_ rbzero.spi_registers.got_new_vinf vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__inv_2
XFILLER_200_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12559_ _05312_ _05314_ _05315_ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__mux2_1
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15278_ _07871_ _07942_ _07963_ vssd1 vssd1 vccd1 vccd1 _07964_ sky130_fd_sc_hd__a21o_1
X_18066_ rbzero.spi_registers.spi_buffer\[9\] rbzero.spi_registers.spi_buffer\[8\]
+ _02227_ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__mux2_1
XFILLER_176_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17017_ rbzero.wall_tracer.trackDistX\[8\] rbzero.wall_tracer.stepDistX\[8\] vssd1
+ vssd1 vccd1 vccd1 _09623_ sky130_fd_sc_hd__or2_1
X_14229_ _06916_ vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__clkbuf_4
XFILLER_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09770_ _02909_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__clkbuf_4
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ rbzero.pov.spi_buffer\[14\] rbzero.pov.ready_buffer\[14\] _02153_ vssd1 vssd1
+ vccd1 vccd1 _02159_ sky130_fd_sc_hd__mux2_1
XFILLER_66_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18899_ _02720_ vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19127__292 clknet_1_0__leaf__02744_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__inv_2
XFILLER_35_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20226_ net286 _01157_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09968_ _03037_ vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__clkbuf_1
X_20157_ net217 _01088_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09899_ _03001_ vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__clkbuf_1
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20088_ clknet_leaf_84_i_clk _01019_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11930_ _04672_ net65 _04704_ _04691_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__a211o_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _04532_ _04635_ _04627_ net14 vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__a31o_1
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13600_ _06354_ _06356_ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__nor2_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10812_ _03589_ _03596_ _03597_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__a21oi_1
XFILLER_72_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _07264_ _07267_ vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__nand2_1
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _04567_ net15 vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__nor2_2
XFILLER_129_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13531_ _05697_ _06055_ vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__and2_1
X_10743_ gpout0.hpos\[0\] _03528_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__or2_1
XFILLER_14_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16250_ _07878_ vssd1 vssd1 vccd1 vccd1 _08862_ sky130_fd_sc_hd__clkbuf_4
XFILLER_159_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13462_ _06215_ _06218_ _06200_ vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__o21a_1
XFILLER_41_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10674_ gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__clkbuf_4
XFILLER_201_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15201_ _07617_ _07646_ _07198_ _07748_ vssd1 vssd1 vccd1 vccd1 _07888_ sky130_fd_sc_hd__or4_1
XFILLER_139_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12413_ _05078_ _05169_ _05072_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__o21a_1
X_16181_ _08788_ _08793_ vssd1 vssd1 vccd1 vccd1 _08794_ sky130_fd_sc_hd__nand2_1
XFILLER_154_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13393_ _05503_ _05987_ vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__or2_1
XFILLER_51_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15132_ _07813_ _07814_ _07815_ _07816_ _07819_ vssd1 vssd1 vccd1 vccd1 _07820_ sky130_fd_sc_hd__o221a_1
XFILLER_127_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12344_ _05039_ _05045_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__or2b_1
XFILLER_114_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19940_ net169 _00871_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[20\] sky130_fd_sc_hd__dfxtp_1
X_15063_ _06759_ _07165_ _06765_ vssd1 vssd1 vccd1 vccd1 _07751_ sky130_fd_sc_hd__o21ai_1
X_12275_ _05031_ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__inv_2
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14014_ _05447_ _06634_ _05322_ vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__a21o_1
XFILLER_107_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11226_ gpout0.vpos\[3\] _03531_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__nor2_1
XFILLER_136_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19871_ clknet_leaf_21_i_clk _00802_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18822_ _04100_ _02634_ vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__and2_1
XFILLER_95_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11157_ rbzero.tex_r1\[45\] _03919_ _03926_ _03673_ vssd1 vssd1 vccd1 vccd1 _03942_
+ sky130_fd_sc_hd__a31o_1
XFILLER_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10108_ _03111_ vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18753_ _02629_ _02413_ _02581_ _02630_ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__a211o_1
X_11088_ rbzero.map_overlay.i_otherx\[2\] vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__inv_2
X_15965_ _08578_ _08579_ _08580_ vssd1 vssd1 vccd1 vccd1 _08581_ sky130_fd_sc_hd__nand3_1
X_17704_ _01971_ _01975_ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__xnor2_1
X_10039_ _03075_ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__clkbuf_1
X_14916_ _07601_ _07603_ _07599_ vssd1 vssd1 vccd1 vccd1 _07604_ sky130_fd_sc_hd__a21oi_1
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18684_ _02575_ _02577_ _02266_ vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__o21a_1
X_15896_ _08513_ _08518_ _08519_ vssd1 vssd1 vccd1 vccd1 _08520_ sky130_fd_sc_hd__nand3b_1
XFILLER_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17635_ _04931_ _01912_ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__xnor2_1
X_14847_ _07532_ _07533_ _07534_ vssd1 vssd1 vccd1 vccd1 _07535_ sky130_fd_sc_hd__o21ba_1
XFILLER_90_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17566_ _01785_ rbzero.wall_tracer.rayAddendY\[7\] vssd1 vssd1 vccd1 vccd1 _01853_
+ sky130_fd_sc_hd__nand2_1
XFILLER_1_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14778_ _07445_ _07462_ vssd1 vssd1 vccd1 vccd1 _07466_ sky130_fd_sc_hd__nor2_1
XFILLER_147_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19305_ rbzero.traced_texa\[-3\] rbzero.texV\[-3\] vssd1 vssd1 vccd1 vccd1 _02794_
+ sky130_fd_sc_hd__nor2_1
X_16517_ _09027_ _09099_ _09126_ vssd1 vssd1 vccd1 vccd1 _09127_ sky130_fd_sc_hd__a21o_1
XFILLER_182_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13729_ _06454_ _06456_ vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18942__126 clknet_1_0__leaf__02725_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__inv_2
X_17497_ _01772_ _01776_ _01787_ _01788_ _03486_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__a311oi_1
XFILLER_17_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16448_ _08922_ _08931_ _08929_ vssd1 vssd1 vccd1 vccd1 _09059_ sky130_fd_sc_hd__a21o_1
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16379_ _08643_ _08081_ vssd1 vssd1 vccd1 vccd1 _08990_ sky130_fd_sc_hd__nor2_1
XFILLER_118_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18118_ rbzero.map_overlay.i_otherx\[2\] _02268_ vssd1 vssd1 vccd1 vccd1 _02269_
+ sky130_fd_sc_hd__or2_1
XFILLER_191_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19098_ clknet_1_0__leaf__02732_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__buf_1
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18049_ _02228_ vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09822_ _02959_ vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__clkbuf_1
X_20011_ clknet_leaf_75_i_clk _00942_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09753_ _02923_ vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19060__232 clknet_1_0__leaf__02737_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__inv_2
XFILLER_23_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10390_ _03259_ vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12060_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__clkinv_2
XFILLER_104_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11011_ _03776_ _03796_ vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__nor2_1
X_20209_ net269 _01140_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12962_ _05689_ _05695_ _05699_ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__nor3_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15750_ _07827_ _08432_ vssd1 vssd1 vccd1 vccd1 _08433_ sky130_fd_sc_hd__xnor2_1
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ _07347_ _07384_ _07388_ vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__a21boi_1
X_11913_ gpout3.clk_div\[1\] _04666_ _04685_ _04687_ vssd1 vssd1 vccd1 vccd1 _04688_
+ sky130_fd_sc_hd__a31o_1
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15681_ _08362_ _08363_ vssd1 vssd1 vccd1 vccd1 _08364_ sky130_fd_sc_hd__and2_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ _05649_ _05648_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__xnor2_2
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _01700_ _01712_ _01701_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__o21ai_1
XFILLER_45_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _07314_ _07309_ vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__or2b_1
X_11844_ _04612_ net67 _04619_ net13 vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a211o_1
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14563_ _07249_ _07250_ vssd1 vssd1 vccd1 vccd1 _07251_ sky130_fd_sc_hd__xnor2_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ rbzero.spi_registers.new_mapd\[4\] rbzero.spi_registers.spi_buffer\[4\] _01663_
+ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__mux2_1
X_11775_ net15 vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__buf_2
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16302_ _08912_ _08913_ vssd1 vssd1 vccd1 vccd1 _08914_ sky130_fd_sc_hd__nand2_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13514_ _06254_ _06269_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__nor2_1
X_10726_ gpout0.hpos\[5\] _03511_ gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1 _03512_
+ sky130_fd_sc_hd__o21a_1
XFILLER_186_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17282_ _01602_ _01607_ vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__nand2_1
X_14494_ _07136_ _07148_ vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__nor2_1
XFILLER_174_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19021_ clknet_1_1__leaf__02732_ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__buf_1
X_16233_ _08760_ _08842_ _08843_ vssd1 vssd1 vccd1 vccd1 _08845_ sky130_fd_sc_hd__and3_1
X_13445_ _06198_ _06201_ vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__xnor2_1
X_10657_ rbzero.map_overlay.i_mapdy\[3\] _03375_ rbzero.map_rom.i_row\[4\] _03451_
+ _03452_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__o221a_1
XFILLER_186_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16164_ _08775_ _08776_ vssd1 vssd1 vccd1 vccd1 _08777_ sky130_fd_sc_hd__xnor2_1
XFILLER_155_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13376_ _06124_ _06127_ _06132_ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10588_ rbzero.wall_tracer.visualWallDist\[7\] rbzero.wall_tracer.visualWallDist\[6\]
+ rbzero.wall_tracer.visualWallDist\[5\] rbzero.wall_tracer.visualWallDist\[4\] vssd1
+ vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__or4_1
XFILLER_127_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15115_ _07336_ _07802_ vssd1 vssd1 vccd1 vccd1 _07803_ sky130_fd_sc_hd__xnor2_4
X_12327_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] vssd1
+ vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__nand2_1
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16095_ _08707_ _08708_ vssd1 vssd1 vccd1 vccd1 _08709_ sky130_fd_sc_hd__xor2_1
XFILLER_114_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15046_ _07094_ _07732_ _07733_ _07093_ vssd1 vssd1 vccd1 vccd1 _07734_ sky130_fd_sc_hd__a22o_1
X_19923_ net152 _00854_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[3\] sky130_fd_sc_hd__dfxtp_1
X_12258_ _05016_ _05014_ _05015_ _05007_ vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__o31ai_1
XFILLER_114_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11209_ _03721_ _03989_ _03993_ _03685_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__a31o_1
XFILLER_96_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19854_ clknet_leaf_23_i_clk _00785_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12189_ rbzero.wall_tracer.state\[1\] _04950_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__nor2_1
X_18805_ _02645_ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__buf_2
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19785_ clknet_leaf_85_i_clk _00716_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[67\]
+ sky130_fd_sc_hd__dfxtp_1
X_16997_ _09601_ _09602_ vssd1 vssd1 vccd1 vccd1 _09603_ sky130_fd_sc_hd__xor2_1
XFILLER_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18736_ rbzero.pov.ready_buffer\[55\] _02413_ _02582_ _02616_ vssd1 vssd1 vccd1 vccd1
+ _02617_ sky130_fd_sc_hd__a211o_1
X_15948_ _08563_ _08564_ _08565_ vssd1 vssd1 vccd1 vccd1 _08566_ sky130_fd_sc_hd__nand3_1
XFILLER_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18667_ rbzero.debug_overlay.playerX\[1\] _02561_ vssd1 vssd1 vccd1 vccd1 _02564_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_64_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15879_ _07826_ _08503_ vssd1 vssd1 vccd1 vccd1 _08505_ sky130_fd_sc_hd__or2_1
XFILLER_110_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17618_ _01899_ vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__clkbuf_1
XFILLER_197_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18598_ _02518_ vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__clkbuf_1
X_17549_ _01836_ _01837_ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__nor2_1
XFILLER_177_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20491_ clknet_leaf_42_i_clk _01422_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_158_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09805_ _02950_ vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__clkbuf_1
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_5_0_i_clk clknet_2_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09736_ _02914_ vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18925__110 clknet_1_0__leaf__02724_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__inv_2
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11560_ _04340_ _04341_ _03659_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__mux2_1
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10511_ _03322_ vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11491_ rbzero.tex_g1\[51\] rbzero.tex_g1\[50\] _04247_ vssd1 vssd1 vccd1 vccd1 _04274_
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13230_ _05950_ _05986_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__xnor2_4
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10442_ _03286_ vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13161_ _05912_ _05917_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__xnor2_1
X_10373_ _03250_ vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12112_ rbzero.debug_overlay.facingY\[0\] rbzero.wall_tracer.rayAddendY\[8\] vssd1
+ vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__nand2_1
XFILLER_163_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13092_ _05836_ _05847_ _05848_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__a21o_1
XFILLER_123_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12043_ _03906_ _03909_ _04790_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__mux2_1
X_16920_ _09520_ _09526_ rbzero.wall_tracer.trackDistX\[7\] _08508_ vssd1 vssd1 vccd1
+ vccd1 _00556_ sky130_fd_sc_hd__o2bb2a_1
X_18971__152 clknet_1_0__leaf__02728_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__inv_2
XFILLER_120_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16851_ _09456_ _09457_ vssd1 vssd1 vccd1 vccd1 _09458_ sky130_fd_sc_hd__nor2_1
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15802_ rbzero.row_render.texu\[4\] _08457_ _08453_ rbzero.wall_tracer.texu\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__a22o_1
X_19570_ clknet_leaf_38_i_clk _00501_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16782_ _09388_ _09389_ vssd1 vssd1 vccd1 vccd1 _09390_ sky130_fd_sc_hd__and2_1
XFILLER_93_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19067__238 clknet_1_1__leaf__02738_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__inv_2
X_13994_ rbzero.wall_tracer.stepDistY\[1\] _06738_ _06718_ vssd1 vssd1 vccd1 vccd1
+ _06739_ sky130_fd_sc_hd__mux2_1
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18521_ _02478_ vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15733_ _08377_ _08415_ vssd1 vssd1 vccd1 vccd1 _08416_ sky130_fd_sc_hd__xnor2_2
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _05669_ _05668_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__and2b_1
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _08202_ _08213_ _08211_ vssd1 vssd1 vccd1 vccd1 _08347_ sky130_fd_sc_hd__a21oi_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _05588_ _05597_ _05632_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__a21o_1
XFILLER_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _01700_ _01701_ vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__and2b_1
XFILLER_33_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14615_ _06919_ _07222_ _07302_ vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__a21bo_1
XFILLER_18_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _04503_ _04552_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__nor2_1
X_15595_ _08276_ _08277_ vssd1 vssd1 vccd1 vccd1 _08279_ sky130_fd_sc_hd__and2_1
XFILLER_18_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _01653_ _01654_ _01652_ vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__a21oi_1
XFILLER_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14546_ _07232_ _07081_ _07233_ vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__o21a_1
XFILLER_92_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11758_ net43 _04516_ _04513_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__and3_1
XFILLER_14_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10709_ _03497_ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__clkbuf_4
X_17265_ rbzero.wall_tracer.trackDistY\[1\] rbzero.wall_tracer.stepDistY\[1\] vssd1
+ vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__or2_1
XFILLER_197_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14477_ _06733_ _07103_ _06752_ _06746_ _06738_ vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__a2111o_2
X_11689_ _04394_ _04469_ _03830_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__mux2_1
XFILLER_146_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16216_ _08601_ _08828_ vssd1 vssd1 vccd1 vccd1 _08829_ sky130_fd_sc_hd__nand2_1
X_13428_ _06182_ _06184_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__and2_1
X_17196_ rbzero.wall_tracer.trackDistY\[-9\] rbzero.wall_tracer.stepDistY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__and2_1
XFILLER_161_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16147_ _08657_ _08729_ _08759_ vssd1 vssd1 vccd1 vccd1 _08760_ sky130_fd_sc_hd__a21o_1
XFILLER_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13359_ _06114_ _06115_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__nand2_1
XFILLER_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16078_ _08690_ _08691_ vssd1 vssd1 vccd1 vccd1 _08692_ sky130_fd_sc_hd__and2b_1
XFILLER_170_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15029_ _07235_ _07052_ vssd1 vssd1 vccd1 vccd1 _07717_ sky130_fd_sc_hd__or2_1
X_19906_ clknet_leaf_25_i_clk _00837_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__04486_ _04486_ vssd1 vssd1 vccd1 vccd1 clknet_0__04486_ sky130_fd_sc_hd__clkbuf_16
X_19837_ clknet_leaf_14_i_clk _00768_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput2 i_debug_vec_overlay vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_6
X_19768_ clknet_leaf_7_i_clk _00699_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18719_ _02603_ _07017_ _02539_ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__mux2_1
X_19699_ clknet_leaf_73_i_clk _00630_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20474_ clknet_leaf_28_i_clk _01405_ vssd1 vssd1 vccd1 vccd1 gpout5.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19172__333 clknet_1_0__leaf__02748_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__inv_2
XFILLER_195_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09719_ _02900_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__clkbuf_4
XFILLER_62_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10991_ rbzero.row_render.size\[7\] rbzero.row_render.size\[6\] vssd1 vssd1 vccd1
+ vccd1 _03777_ sky130_fd_sc_hd__xnor2_1
XFILLER_55_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12730_ _05475_ _05486_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__xnor2_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _05378_ _05384_ _05329_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__a21o_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _04911_ _05086_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__mux2_1
X_11612_ _04393_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__inv_2
XFILLER_187_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ _07790_ _07844_ _07966_ _07964_ vssd1 vssd1 vccd1 vccd1 _08065_ sky130_fd_sc_hd__o31ai_2
X_12592_ _05311_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__clkbuf_4
XFILLER_129_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11543_ rbzero.tex_b0\[49\] rbzero.tex_b0\[48\] _03732_ vssd1 vssd1 vccd1 vccd1 _04325_
+ sky130_fd_sc_hd__mux2_1
X_14331_ _03492_ _07018_ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__nand2_1
XFILLER_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17050_ _09280_ _09634_ _09633_ vssd1 vssd1 vccd1 vccd1 _09655_ sky130_fd_sc_hd__o21ba_1
X_14262_ rbzero.wall_tracer.state\[13\] rbzero.wall_tracer.stepDistY\[-6\] rbzero.wall_tracer.state\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__a21o_1
X_11474_ rbzero.tex_g1\[13\] rbzero.tex_g1\[12\] _03618_ vssd1 vssd1 vccd1 vccd1 _04257_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16001_ _08613_ _08614_ vssd1 vssd1 vccd1 vccd1 _08615_ sky130_fd_sc_hd__xnor2_1
X_13213_ _05927_ _05969_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__xnor2_1
XFILLER_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10425_ _03277_ vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14193_ rbzero.wall_tracer.visualWallDist\[-7\] _06880_ rbzero.wall_tracer.state\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__mux2_1
XFILLER_164_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13144_ _05852_ _05855_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__xor2_2
XFILLER_100_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10356_ _03241_ vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13075_ _05825_ _05829_ _05831_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__o21ai_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17952_ _02176_ vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__clkbuf_1
X_10287_ _03205_ vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16903_ _09320_ _09399_ _09509_ vssd1 vssd1 vccd1 vccd1 _09510_ sky130_fd_sc_hd__a21oi_1
X_12026_ net47 net48 _03910_ net69 _04790_ _04792_ vssd1 vssd1 vccd1 vccd1 _04799_
+ sky130_fd_sc_hd__mux4_1
XFILLER_39_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17883_ _02137_ _02103_ _02138_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__and3b_1
XFILLER_93_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19622_ clknet_leaf_48_i_clk _00553_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16834_ _09439_ _09440_ vssd1 vssd1 vccd1 vccd1 _09441_ sky130_fd_sc_hd__nand2_1
XFILLER_120_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19553_ clknet_leaf_34_i_clk _00484_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[3\] sky130_fd_sc_hd__dfxtp_1
X_16765_ _09356_ _09277_ _09371_ vssd1 vssd1 vccd1 vccd1 _09373_ sky130_fd_sc_hd__nand3_1
XFILLER_81_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13977_ _06721_ _06690_ _06708_ _06723_ _06664_ _05310_ vssd1 vssd1 vccd1 vccd1 _06724_
+ sky130_fd_sc_hd__mux4_1
XFILLER_111_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18504_ _02469_ vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15716_ _06860_ _08397_ _07162_ _08398_ _04841_ vssd1 vssd1 vccd1 vccd1 _08399_ sky130_fd_sc_hd__o221a_1
XFILLER_111_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12928_ _05682_ _05683_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__or2b_1
X_19484_ clknet_leaf_57_i_clk _00430_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
X_16696_ _09191_ _09193_ vssd1 vssd1 vccd1 vccd1 _09305_ sky130_fd_sc_hd__or2_1
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15647_ _08328_ _08329_ vssd1 vssd1 vccd1 vccd1 _08330_ sky130_fd_sc_hd__or2_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _05469_ _05615_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__nand2_2
XFILLER_61_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18366_ rbzero.pov.spi_counter\[2\] _02417_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__and2_1
XFILLER_159_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15578_ _08259_ _08261_ vssd1 vssd1 vccd1 vccd1 _08262_ sky130_fd_sc_hd__nand2_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17317_ rbzero.wall_tracer.trackDistY\[8\] rbzero.wall_tracer.stepDistY\[8\] vssd1
+ vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__nand2_1
XFILLER_119_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14529_ _07196_ _07214_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__nand2_1
X_18297_ rbzero.spi_registers.spi_buffer\[2\] rbzero.spi_registers.new_leak\[2\] _02379_
+ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__mux2_1
XFILLER_175_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17248_ _01578_ _01579_ _01580_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__a21o_1
XFILLER_174_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18978__158 clknet_1_1__leaf__02729_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__inv_2
XFILLER_127_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17179_ rbzero.wall_tracer.state\[1\] _03493_ _01521_ vssd1 vssd1 vccd1 vccd1 _01522_
+ sky130_fd_sc_hd__o21a_2
XFILLER_127_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20190_ net250 _01121_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_40 net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_51 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_62 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20457_ net137 _01388_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[48\] sky130_fd_sc_hd__dfxtp_1
X_10210_ rbzero.tex_g0\[29\] rbzero.tex_g0\[28\] _03155_ vssd1 vssd1 vccd1 vccd1 _03165_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11190_ rbzero.tex_r1\[8\] _03920_ _03925_ _03973_ _03974_ vssd1 vssd1 vccd1 vccd1
+ _03975_ sky130_fd_sc_hd__a311o_1
X_20388_ net448 _01319_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10141_ _03128_ vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10072_ _03092_ vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13900_ _06619_ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__inv_2
XFILLER_101_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14880_ _07545_ _07567_ vssd1 vssd1 vccd1 vccd1 _07568_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_2_0_i_clk clknet_1_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_130_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13831_ _05324_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__buf_2
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16550_ _09158_ _09159_ vssd1 vssd1 vccd1 vccd1 _09160_ sky130_fd_sc_hd__xnor2_1
XFILLER_56_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10974_ rbzero.tex_r0\[50\] _03700_ _03659_ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__a21o_1
X_13762_ _05551_ _06230_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__nor2_1
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15501_ _08065_ _08169_ _08184_ vssd1 vssd1 vccd1 vccd1 _08185_ sky130_fd_sc_hd__a21o_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12713_ _05355_ _05469_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__xor2_1
X_16481_ _09075_ _08967_ vssd1 vssd1 vccd1 vccd1 _09091_ sky130_fd_sc_hd__and2b_1
X_13693_ _06446_ _06449_ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__nor2_1
XFILLER_16_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18220_ _04827_ vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__buf_4
X_15432_ _08007_ _08010_ vssd1 vssd1 vccd1 vccd1 _08117_ sky130_fd_sc_hd__or2b_1
X_12644_ _05347_ _05400_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__nor2_1
XFILLER_62_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19179__339 clknet_1_1__leaf__02749_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__inv_2
XFILLER_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18151_ rbzero.map_overlay.i_mapdx\[0\] _02292_ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__or2_1
XFILLER_50_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12575_ _05330_ _05331_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__and2_1
X_15363_ _07927_ vssd1 vssd1 vccd1 vccd1 _08049_ sky130_fd_sc_hd__inv_2
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17102_ _09615_ _09619_ _09613_ vssd1 vssd1 vccd1 vccd1 _09707_ sky130_fd_sc_hd__a21o_1
XFILLER_184_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14314_ _06849_ _04898_ vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__nor2_1
XFILLER_141_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18082_ rbzero.spi_registers.mosi _02107_ _02245_ vssd1 vssd1 vccd1 vccd1 _02246_
+ sky130_fd_sc_hd__mux2_1
X_11526_ _04235_ _04308_ _03830_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__mux2_1
X_15294_ _07078_ _07273_ _07092_ _07039_ vssd1 vssd1 vccd1 vccd1 _07980_ sky130_fd_sc_hd__o22a_1
XFILLER_8_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17033_ _09007_ _09035_ _09036_ _09009_ vssd1 vssd1 vccd1 vccd1 _09638_ sky130_fd_sc_hd__o22ai_1
XFILLER_8_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11457_ rbzero.tex_g1\[19\] rbzero.tex_g1\[18\] _03617_ vssd1 vssd1 vccd1 vccd1 _04240_
+ sky130_fd_sc_hd__mux2_1
X_14245_ _06932_ vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__clkbuf_4
XFILLER_125_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10408_ _03268_ vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__clkbuf_1
X_14176_ _06860_ rbzero.wall_tracer.stepDistY\[-11\] _06863_ _04840_ vssd1 vssd1 vccd1
+ vccd1 _06864_ sky130_fd_sc_hd__o211a_1
XFILLER_194_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11388_ rbzero.tex_g0\[1\] rbzero.tex_g0\[0\] _03615_ vssd1 vssd1 vccd1 vccd1 _04172_
+ sky130_fd_sc_hd__mux2_1
XFILLER_178_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ rbzero.tex_b1\[31\] rbzero.tex_b1\[32\] _03232_ vssd1 vssd1 vccd1 vccd1 _03233_
+ sky130_fd_sc_hd__mux2_1
X_13127_ _05882_ _05883_ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__and2_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17935_ _02167_ vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__clkbuf_1
X_13058_ _05804_ _05808_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__or2_1
XFILLER_79_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12009_ _04779_ net67 _04781_ net37 vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__a211o_1
XFILLER_66_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17866_ rbzero.spi_registers.spi_counter\[1\] _02102_ _02103_ _02125_ vssd1 vssd1
+ vccd1 vccd1 _00643_ sky130_fd_sc_hd__o211a_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16817_ _09353_ _09322_ vssd1 vssd1 vccd1 vccd1 _09424_ sky130_fd_sc_hd__or2b_1
X_19605_ clknet_leaf_63_i_clk _00536_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_17797_ _02000_ rbzero.wall_tracer.rayAddendX\[7\] vssd1 vssd1 vccd1 vccd1 _02062_
+ sky130_fd_sc_hd__nand2_1
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19536_ clknet_leaf_38_i_clk _00007_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_16748_ _09269_ _09275_ vssd1 vssd1 vccd1 vccd1 _09356_ sky130_fd_sc_hd__nand2_1
XFILLER_62_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19467_ clknet_leaf_61_i_clk _00413_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16679_ _09286_ _09287_ vssd1 vssd1 vccd1 vccd1 _09288_ sky130_fd_sc_hd__nor2_1
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19398_ rbzero.traced_texVinit\[4\] _02868_ _08052_ _01745_ vssd1 vssd1 vccd1 vccd1
+ _01432_ sky130_fd_sc_hd__a22o_1
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18349_ rbzero.spi_registers.got_new_vinf _02323_ _02283_ _02408_ vssd1 vssd1 vccd1
+ vccd1 _00842_ sky130_fd_sc_hd__a31o_1
XFILLER_147_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20311_ net371 _01242_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_6_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_190_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20242_ net302 _01173_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20173_ net233 _01104_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[20\] sky130_fd_sc_hd__dfxtp_1
X_09984_ rbzero.tex_r0\[8\] rbzero.tex_r0\[7\] _03039_ vssd1 vssd1 vccd1 vccd1 _03046_
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10690_ rbzero.wall_tracer.state\[0\] vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__inv_2
XFILLER_179_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12360_ rbzero.wall_tracer.visualWallDist\[-10\] rbzero.wall_tracer.rayAddendY\[-2\]
+ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__mux2_1
XFILLER_194_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11311_ rbzero.debug_overlay.facingY\[10\] _04078_ _04088_ _04095_ vssd1 vssd1 vccd1
+ vccd1 _04096_ sky130_fd_sc_hd__a211o_1
XFILLER_126_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20509_ clknet_leaf_30_i_clk _01440_ vssd1 vssd1 vccd1 vccd1 gpout0.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12291_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] _05047_
+ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__a21o_1
XFILLER_10_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14030_ _05322_ _06724_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__nand2_1
X_11242_ _04024_ _04026_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__and2b_1
XFILLER_10_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11173_ _03685_ _03929_ _03939_ _03957_ _03719_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__o311a_1
XFILLER_164_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10124_ rbzero.tex_g1\[5\] rbzero.tex_g1\[6\] _03117_ vssd1 vssd1 vccd1 vccd1 _03120_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15981_ _08592_ _08593_ _08594_ _08589_ vssd1 vssd1 vccd1 vccd1 _08595_ sky130_fd_sc_hd__o211a_1
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17720_ _04100_ rbzero.debug_overlay.vplaneX\[-9\] _01979_ vssd1 vssd1 vccd1 vccd1
+ _01991_ sky130_fd_sc_hd__a21oi_1
X_14932_ _07577_ _07618_ _07619_ vssd1 vssd1 vccd1 vccd1 _07620_ sky130_fd_sc_hd__o21a_1
X_10055_ _03083_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17651_ rbzero.debug_overlay.vplaneX\[-6\] rbzero.wall_tracer.rayAddendX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__nand2_1
XFILLER_75_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14863_ _07502_ _07510_ vssd1 vssd1 vccd1 vccd1 _07551_ sky130_fd_sc_hd__xor2_1
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16602_ _09109_ _09125_ _09123_ vssd1 vssd1 vccd1 vccd1 _09211_ sky130_fd_sc_hd__a21o_1
XFILLER_21_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13814_ _06227_ _06570_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__xor2_1
XFILLER_91_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17582_ _01853_ _01858_ _01867_ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__a21oi_1
X_14794_ _07101_ _06969_ vssd1 vssd1 vccd1 vccd1 _07482_ sky130_fd_sc_hd__nor2_1
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19321_ _02800_ _02802_ _02801_ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__a21boi_1
XFILLER_189_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16533_ _08108_ _09142_ vssd1 vssd1 vccd1 vccd1 _09143_ sky130_fd_sc_hd__nor2_1
X_13745_ _06500_ _06501_ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__and2_1
XFILLER_91_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10957_ _03611_ _03742_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__or2_1
XFILLER_44_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16464_ _08844_ _09074_ vssd1 vssd1 vccd1 vccd1 _09075_ sky130_fd_sc_hd__xnor2_2
XFILLER_149_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13676_ _06432_ _06431_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__nor2_1
X_10888_ _03673_ vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__buf_6
XFILLER_188_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18203_ _02322_ vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__clkbuf_1
X_15415_ _07865_ _07857_ vssd1 vssd1 vccd1 vccd1 _08100_ sky130_fd_sc_hd__nor2_1
X_12627_ _05217_ _05305_ _05302_ _05306_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__or4_1
X_16395_ _08891_ _08903_ _08901_ vssd1 vssd1 vccd1 vccd1 _09006_ sky130_fd_sc_hd__a21o_1
XFILLER_129_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18134_ rbzero.spi_registers.new_other\[4\] _02264_ _02277_ _02275_ vssd1 vssd1 vccd1
+ vccd1 _00759_ sky130_fd_sc_hd__o211a_1
XFILLER_89_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15346_ _08006_ _08031_ vssd1 vssd1 vccd1 vccd1 _08032_ sky130_fd_sc_hd__xnor2_2
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12558_ _05304_ _05299_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__xnor2_4
XFILLER_8_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11509_ _04290_ _04291_ _03920_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__mux2_1
X_18065_ _02236_ vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__clkbuf_1
X_15277_ _07958_ _07962_ vssd1 vssd1 vccd1 vccd1 _07963_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12489_ _05224_ _05226_ _05232_ _05245_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__or4_2
XFILLER_176_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17016_ _09615_ _09619_ _09621_ vssd1 vssd1 vccd1 vccd1 _09622_ sky130_fd_sc_hd__o21ai_2
XFILLER_176_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14228_ _06906_ _06911_ _06913_ _06915_ vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_171_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14159_ _03458_ _06847_ _06848_ _00016_ vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__o22a_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17918_ _02158_ vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__clkbuf_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18898_ _02334_ _02718_ _02719_ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__and3_1
XFILLER_39_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17849_ rbzero.spi_registers.spi_cmd\[3\] rbzero.spi_registers.spi_cmd\[2\] vssd1
+ vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__nor2_1
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19519_ clknet_leaf_49_i_clk _00465_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20225_ net285 _01156_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20156_ net216 _01087_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09967_ rbzero.tex_r0\[16\] rbzero.tex_r0\[15\] _03028_ vssd1 vssd1 vccd1 vccd1 _03037_
+ sky130_fd_sc_hd__mux2_1
XFILLER_103_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20087_ clknet_leaf_84_i_clk _01018_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09898_ rbzero.tex_r0\[49\] rbzero.tex_r0\[48\] _02995_ vssd1 vssd1 vccd1 vccd1 _03001_
+ sky130_fd_sc_hd__mux2_1
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ net44 _04625_ _04623_ _04634_ _04635_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__a32o_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _03586_ _03588_ _03585_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__a21oi_1
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11791_ _04567_ net15 vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__and2_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13530_ _06246_ _06248_ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__xnor2_1
XFILLER_40_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10742_ _03526_ _03527_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__or2_1
XFILLER_158_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13461_ _06217_ vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__inv_2
X_10673_ _03461_ _02901_ _03465_ _03467_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__o31a_1
XFILLER_185_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15200_ _07100_ _07137_ vssd1 vssd1 vccd1 vccd1 _07887_ sky130_fd_sc_hd__or2_1
XFILLER_22_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12412_ rbzero.wall_tracer.visualWallDist\[9\] _03480_ vssd1 vssd1 vccd1 vccd1 _05169_
+ sky130_fd_sc_hd__nor2_1
XFILLER_167_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16180_ _08791_ _08792_ vssd1 vssd1 vccd1 vccd1 _08793_ sky130_fd_sc_hd__xor2_1
XFILLER_139_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13392_ _06001_ _05992_ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__nor2_1
XFILLER_12_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15131_ _07817_ _07818_ _07815_ _07816_ vssd1 vssd1 vccd1 vccd1 _07819_ sky130_fd_sc_hd__a22o_1
XFILLER_182_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12343_ _05038_ _05044_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__nor2_1
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12274_ rbzero.debug_overlay.facingX\[-4\] rbzero.wall_tracer.rayAddendX\[4\] vssd1
+ vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__nand2_1
XFILLER_5_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15062_ _06759_ _06764_ _07165_ vssd1 vssd1 vccd1 vccd1 _07750_ sky130_fd_sc_hd__or3_1
XFILLER_154_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11225_ _04008_ _04009_ _03902_ _03461_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__o211a_1
X_14013_ _06675_ _06730_ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__nor2_1
XFILLER_175_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19870_ clknet_leaf_3_i_clk _00801_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_done
+ sky130_fd_sc_hd__dfxtp_1
X_11156_ rbzero.tex_r1\[47\] _03664_ _03940_ _03677_ vssd1 vssd1 vccd1 vccd1 _03941_
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18821_ rbzero.pov.ready_buffer\[14\] _02663_ _02671_ _02672_ vssd1 vssd1 vccd1 vccd1
+ _01051_ sky130_fd_sc_hd__o211a_1
XFILLER_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10107_ rbzero.tex_g1\[13\] rbzero.tex_g1\[14\] _03106_ vssd1 vssd1 vccd1 vccd1 _03111_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18752_ rbzero.debug_overlay.playerY\[5\] rbzero.debug_overlay.playerY\[4\] _02619_
+ _02539_ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__o31a_1
X_11087_ rbzero.map_overlay.i_othery\[3\] vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__inv_2
X_15964_ _08570_ _08572_ _08571_ vssd1 vssd1 vccd1 vccd1 _08580_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17703_ _01973_ _01974_ vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__or2_1
X_10038_ rbzero.tex_g1\[46\] rbzero.tex_g1\[47\] _03073_ vssd1 vssd1 vccd1 vccd1 _03075_
+ sky130_fd_sc_hd__mux2_1
X_14915_ _07583_ _07602_ vssd1 vssd1 vccd1 vccd1 _07603_ sky130_fd_sc_hd__nor2_1
X_18683_ rbzero.pov.ready_buffer\[72\] _02540_ _02543_ _02576_ vssd1 vssd1 vccd1 vccd1
+ _02577_ sky130_fd_sc_hd__o211a_1
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15895_ rbzero.wall_tracer.trackDistX\[-10\] rbzero.wall_tracer.stepDistX\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _08519_ sky130_fd_sc_hd__nand2_1
XFILLER_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17634_ rbzero.map_rom.i_row\[4\] _04923_ _04943_ vssd1 vssd1 vccd1 vccd1 _01912_
+ sky130_fd_sc_hd__a21oi_1
X_14846_ _07119_ _06917_ _06978_ _07005_ vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__nor4_1
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17565_ _08458_ _01843_ _01844_ _01852_ vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__a31o_1
XFILLER_91_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14777_ _07443_ _07464_ vssd1 vssd1 vccd1 vccd1 _07465_ sky130_fd_sc_hd__nor2_1
X_11989_ net40 _04730_ _04732_ _03537_ _04762_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__a221o_1
XFILLER_90_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19304_ rbzero.texV\[-4\] _02675_ _02709_ _02793_ vssd1 vssd1 vccd1 vccd1 _01413_
+ sky130_fd_sc_hd__a22o_1
X_16516_ _09109_ _09125_ vssd1 vssd1 vccd1 vccd1 _09126_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13728_ _06483_ _06484_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__xnor2_1
XFILLER_56_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17496_ _01772_ _01776_ _01787_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16447_ _09045_ _09057_ vssd1 vssd1 vccd1 vccd1 _09058_ sky130_fd_sc_hd__xnor2_2
X_13659_ _06406_ _06415_ _06413_ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__a21o_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_158_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16378_ _08865_ _08987_ _08988_ vssd1 vssd1 vccd1 vccd1 _08989_ sky130_fd_sc_hd__a21bo_1
XFILLER_191_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18117_ rbzero.spi_registers.got_new_other _02262_ vssd1 vssd1 vccd1 vccd1 _02268_
+ sky130_fd_sc_hd__and2_1
X_15329_ _04832_ _08013_ _08014_ _07162_ vssd1 vssd1 vccd1 vccd1 _08015_ sky130_fd_sc_hd__a31o_1
XFILLER_145_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18048_ rbzero.spi_registers.spi_buffer\[0\] rbzero.spi_registers.mosi _02227_ vssd1
+ vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__mux2_1
XFILLER_132_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_86_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_126_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20010_ clknet_leaf_75_i_clk _00941_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09821_ rbzero.tex_r1\[19\] rbzero.tex_r1\[20\] _02954_ vssd1 vssd1 vccd1 vccd1 _02959_
+ sky130_fd_sc_hd__mux2_1
XFILLER_141_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19999_ clknet_leaf_93_i_clk _00930_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09752_ rbzero.tex_r1\[52\] rbzero.tex_r1\[53\] _02921_ vssd1 vssd1 vccd1 vccd1 _02923_
+ sky130_fd_sc_hd__mux2_1
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_81_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_39_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_149_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_1_0_i_clk clknet_2_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_183_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11010_ rbzero.row_render.size\[8\] rbzero.row_render.size\[7\] _03775_ vssd1 vssd1
+ vccd1 vccd1 _03796_ sky130_fd_sc_hd__nor3_1
X_20208_ net268 _01139_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20139_ clknet_leaf_0_i_clk _01070_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_done sky130_fd_sc_hd__dfxtp_1
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12961_ _05716_ _05717_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__xor2_1
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _07385_ _07387_ vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__nand2_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11912_ net46 _04665_ _04685_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__and3_1
X_15680_ _08224_ _08361_ vssd1 vssd1 vccd1 vccd1 _08363_ sky130_fd_sc_hd__or2_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _05493_ _05550_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__or2_1
XFILLER_18_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _06876_ _07014_ _07061_ _07060_ vssd1 vssd1 vccd1 vccd1 _07319_ sky130_fd_sc_hd__a31o_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _04612_ _03913_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__nor2_1
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17350_ _01667_ vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__clkbuf_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _07007_ _07052_ vssd1 vssd1 vccd1 vccd1 _07250_ sky130_fd_sc_hd__or2_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _04498_ _04526_ _04550_ _04551_ vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__o31a_2
XFILLER_199_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _08245_ _08260_ _08018_ _08247_ vssd1 vssd1 vccd1 vccd1 _08913_ sky130_fd_sc_hd__o22ai_1
XFILLER_158_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13513_ _06254_ _06269_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__xor2_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ gpout0.hpos\[4\] _03503_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__or2_1
X_17281_ rbzero.wall_tracer.trackDistY\[3\] rbzero.wall_tracer.stepDistY\[3\] vssd1
+ vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__or2_1
XFILLER_201_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14493_ _07155_ _07180_ vssd1 vssd1 vccd1 vccd1 _07181_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16232_ _08760_ _08842_ _08843_ vssd1 vssd1 vccd1 vccd1 _08844_ sky130_fd_sc_hd__a21oi_2
XFILLER_158_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13444_ _06082_ _06110_ _06199_ _06200_ vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__o31a_1
XFILLER_186_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10656_ rbzero.map_overlay.i_mapdy\[0\] _03390_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__xnor2_1
XFILLER_167_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16163_ _08108_ _08252_ vssd1 vssd1 vccd1 vccd1 _08776_ sky130_fd_sc_hd__or2_1
X_13375_ _06127_ _06131_ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__nor2_1
X_10587_ _03372_ _03377_ _03380_ _03382_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__or4_1
XFILLER_155_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15114_ _07799_ _07801_ vssd1 vssd1 vccd1 vccd1 _07802_ sky130_fd_sc_hd__xor2_4
XFILLER_154_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12326_ _05034_ _05037_ _05046_ _05050_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__a31o_1
X_16094_ _08320_ _08423_ _08421_ vssd1 vssd1 vccd1 vccd1 _08708_ sky130_fd_sc_hd__a21oi_1
XFILLER_108_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15045_ _06970_ _07141_ vssd1 vssd1 vccd1 vccd1 _07733_ sky130_fd_sc_hd__nor2_1
X_19922_ net151 _00853_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12257_ _05014_ _05015_ _05016_ vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__o21a_1
X_11208_ rbzero.tex_r1\[16\] _03920_ _03925_ _03991_ _03992_ vssd1 vssd1 vccd1 vccd1
+ _03993_ sky130_fd_sc_hd__a311o_1
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19237__12 clknet_1_0__leaf__02754_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__inv_2
XFILLER_122_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19853_ clknet_leaf_21_i_clk _00784_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12188_ _04949_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__clkbuf_4
XFILLER_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18804_ rbzero.pov.ready_buffer\[29\] _02644_ _02662_ _02651_ vssd1 vssd1 vccd1 vccd1
+ _01044_ sky130_fd_sc_hd__a211o_1
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11139_ rbzero.tex_r1\[51\] _03618_ _03923_ _03917_ vssd1 vssd1 vccd1 vccd1 _03924_
+ sky130_fd_sc_hd__o211a_1
XFILLER_23_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16996_ _09464_ _09502_ _09501_ vssd1 vssd1 vccd1 vccd1 _09602_ sky130_fd_sc_hd__o21ba_1
X_19784_ clknet_leaf_82_i_clk _00715_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19252__26 clknet_1_1__leaf__02755_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__inv_2
XFILLER_23_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18735_ _02614_ _02615_ _02412_ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__a21oi_1
XFILLER_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15947_ _08555_ _08557_ _08556_ vssd1 vssd1 vccd1 vccd1 _08565_ sky130_fd_sc_hd__o21bai_1
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18666_ rbzero.debug_overlay.playerX\[0\] _02534_ _02563_ _02559_ vssd1 vssd1 vccd1
+ vccd1 _01005_ sky130_fd_sc_hd__a211o_1
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15878_ _07826_ _08503_ vssd1 vssd1 vccd1 vccd1 _08504_ sky130_fd_sc_hd__nand2_1
XFILLER_92_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17617_ _01898_ _03358_ _05009_ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__mux2_1
X_14829_ _07499_ _07516_ vssd1 vssd1 vccd1 vccd1 _07517_ sky130_fd_sc_hd__xor2_1
X_19044__217 clknet_1_0__leaf__02736_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__inv_2
X_18597_ rbzero.pov.spi_buffer\[66\] rbzero.pov.spi_buffer\[67\] _02510_ vssd1 vssd1
+ vccd1 vccd1 _02518_ sky130_fd_sc_hd__mux2_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17548_ _01818_ _01834_ _01835_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__nor3_1
XFILLER_189_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17479_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__nand2_1
XFILLER_177_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20490_ clknet_leaf_42_i_clk _01421_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19090__259 clknet_1_0__leaf__02740_ vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__inv_2
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09804_ rbzero.tex_r1\[27\] rbzero.tex_r1\[28\] _02943_ vssd1 vssd1 vccd1 vccd1 _02950_
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18436__76 clknet_1_1__leaf__02438_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__inv_2
XFILLER_189_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09735_ rbzero.tex_r1\[60\] rbzero.tex_r1\[61\] _02910_ vssd1 vssd1 vccd1 vccd1 _02914_
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10510_ rbzero.tex_b0\[14\] rbzero.tex_b0\[13\] _03313_ vssd1 vssd1 vccd1 vccd1 _03322_
+ sky130_fd_sc_hd__mux2_1
X_11490_ _03721_ _04260_ _04264_ _04272_ _03685_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__o311a_1
XFILLER_156_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10441_ rbzero.tex_b0\[47\] rbzero.tex_b0\[46\] _03280_ vssd1 vssd1 vccd1 vccd1 _03286_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10372_ rbzero.tex_b1\[15\] rbzero.tex_b1\[16\] _03243_ vssd1 vssd1 vccd1 vccd1 _03250_
+ sky130_fd_sc_hd__mux2_1
X_13160_ _05913_ _05916_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12111_ _04865_ _04869_ _04872_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__a21oi_2
X_13091_ _05801_ _05835_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__and2_1
XFILLER_123_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12042_ _04814_ _04787_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__or2b_1
XFILLER_123_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16850_ _09454_ _09455_ vssd1 vssd1 vccd1 vccd1 _09457_ sky130_fd_sc_hd__and2_1
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15801_ rbzero.row_render.texu\[3\] _08457_ _08453_ rbzero.wall_tracer.texu\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__a22o_1
XFILLER_59_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16781_ _09386_ _09387_ vssd1 vssd1 vccd1 vccd1 _09389_ sky130_fd_sc_hd__nand2_1
XFILLER_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13993_ _05320_ _06673_ _06736_ _05390_ _06737_ vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__o221ai_4
XFILLER_92_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18520_ rbzero.pov.spi_buffer\[29\] rbzero.pov.spi_buffer\[30\] _02477_ vssd1 vssd1
+ vccd1 vccd1 _02478_ sky130_fd_sc_hd__mux2_1
X_15732_ _08413_ _08414_ vssd1 vssd1 vccd1 vccd1 _08415_ sky130_fd_sc_hd__and2b_1
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ _05671_ _05672_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__xnor2_1
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15663_ _08336_ _08345_ vssd1 vssd1 vccd1 vccd1 _08346_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12875_ _05589_ _05596_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__and2b_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17402_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.wall_tracer.rayAddendY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__nand2_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _06908_ _06917_ _07220_ vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__or3_1
X_18382_ clknet_1_1__leaf__02433_ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__buf_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ net17 _04602_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__nand2_1
X_15594_ _08276_ _08277_ vssd1 vssd1 vccd1 vccd1 _08278_ sky130_fd_sc_hd__nor2_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17333_ _01652_ _01653_ _01654_ vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__and3_1
XFILLER_18_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14545_ _06900_ _06940_ _06968_ _06970_ vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__or4_1
XFILLER_53_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ net48 _04515_ _04516_ net47 vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__a22o_1
XFILLER_186_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10708_ _03484_ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__buf_6
X_17264_ rbzero.wall_tracer.trackDistY\[1\] rbzero.wall_tracer.stepDistY\[1\] vssd1
+ vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__nand2_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14476_ _06733_ _07103_ _06746_ _06738_ vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__a211oi_1
X_11688_ _03764_ _04396_ _04398_ _04433_ _04468_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__o32a_1
XFILLER_201_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16215_ _08826_ _08827_ vssd1 vssd1 vccd1 vccd1 _08828_ sky130_fd_sc_hd__xor2_1
X_13427_ _06181_ _06176_ _06180_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__nand3_1
X_10639_ rbzero.map_overlay.i_othery\[3\] rbzero.map_rom.a6 vssd1 vssd1 vccd1 vccd1
+ _03435_ sky130_fd_sc_hd__xor2_1
X_17195_ rbzero.wall_tracer.trackDistY\[-9\] rbzero.wall_tracer.stepDistY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__nor2_1
X_16146_ _08741_ _08758_ vssd1 vssd1 vccd1 vccd1 _08759_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13358_ _06096_ _06113_ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__or2_1
XFILLER_182_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12309_ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__inv_2
XFILLER_170_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16077_ _08687_ _08689_ vssd1 vssd1 vccd1 vccd1 _08691_ sky130_fd_sc_hd__nand2_1
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13289_ _06020_ _06045_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__xor2_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15028_ _07714_ _07715_ vssd1 vssd1 vccd1 vccd1 _07716_ sky130_fd_sc_hd__nand2_1
X_19905_ clknet_leaf_23_i_clk _00836_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19836_ clknet_leaf_14_i_clk _00767_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdy\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19767_ clknet_leaf_7_i_clk _00698_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_16979_ _09583_ _09584_ vssd1 vssd1 vccd1 vccd1 _09585_ sky130_fd_sc_hd__xnor2_1
Xinput3 i_gpout0_sel[0] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_6
XFILLER_49_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18718_ rbzero.pov.ready_buffer\[51\] vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__inv_2
XFILLER_25_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19698_ clknet_leaf_73_i_clk _00629_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18649_ rbzero.pov.ready_buffer\[64\] _06963_ _02539_ vssd1 vssd1 vccd1 vccd1 _02551_
+ sky130_fd_sc_hd__mux2_1
XFILLER_149_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20473_ clknet_leaf_28_i_clk _01404_ vssd1 vssd1 vccd1 vccd1 gpout5.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18955__137 clknet_1_0__leaf__02727_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__inv_2
XFILLER_160_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09718_ gpout0.hpos\[7\] vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__buf_4
X_10990_ rbzero.row_render.size\[7\] _03775_ rbzero.row_render.size\[8\] vssd1 vssd1
+ vccd1 vccd1 _03776_ sky130_fd_sc_hd__o21a_1
XFILLER_167_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _05414_ _05363_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__or2_2
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _03522_ _04392_ _03912_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__o21ai_4
XFILLER_42_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12591_ _05180_ _05181_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__nand2_1
XFILLER_169_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14330_ rbzero.debug_overlay.playerY\[-2\] _07017_ _04928_ vssd1 vssd1 vccd1 vccd1
+ _07018_ sky130_fd_sc_hd__mux2_1
XFILLER_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11542_ rbzero.tex_b0\[51\] rbzero.tex_b0\[50\] _03732_ vssd1 vssd1 vccd1 vccd1 _04324_
+ sky130_fd_sc_hd__mux2_1
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14261_ _04947_ _06945_ _06947_ _06948_ vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_183_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11473_ _03648_ _04246_ _04255_ _03688_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__o211a_1
XFILLER_7_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16000_ _07269_ _08316_ vssd1 vssd1 vccd1 vccd1 _08614_ sky130_fd_sc_hd__and2_1
XFILLER_100_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13212_ _05961_ _05968_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10424_ rbzero.tex_b0\[55\] rbzero.tex_b0\[54\] _03269_ vssd1 vssd1 vccd1 vccd1 _03277_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14192_ rbzero.debug_overlay.playerY\[-7\] _06879_ _04927_ vssd1 vssd1 vccd1 vccd1
+ _06880_ sky130_fd_sc_hd__mux2_1
XFILLER_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13143_ _05856_ _05899_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__xnor2_1
X_10355_ rbzero.tex_b1\[23\] rbzero.tex_b1\[24\] _03232_ vssd1 vssd1 vccd1 vccd1 _03241_
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ rbzero.tex_b1\[56\] rbzero.tex_b1\[57\] _03199_ vssd1 vssd1 vccd1 vccd1 _03205_
+ sky130_fd_sc_hd__mux2_1
XFILLER_174_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13074_ _05795_ _05830_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__nor2_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17951_ rbzero.pov.spi_buffer\[29\] rbzero.pov.ready_buffer\[29\] _02175_ vssd1 vssd1
+ vccd1 vccd1 _02176_ sky130_fd_sc_hd__mux2_1
XFILLER_78_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16902_ _09396_ _09398_ vssd1 vssd1 vccd1 vccd1 _09509_ sky130_fd_sc_hd__nor2_1
X_12025_ net36 vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__inv_2
X_17882_ rbzero.spi_registers.spi_counter\[5\] _02136_ vssd1 vssd1 vccd1 vccd1 _02138_
+ sky130_fd_sc_hd__or2_1
XFILLER_39_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19621_ clknet_leaf_47_i_clk _00552_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16833_ _08643_ _08317_ vssd1 vssd1 vccd1 vccd1 _09440_ sky130_fd_sc_hd__and2_1
XFILLER_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16764_ _09356_ _09277_ _09371_ vssd1 vssd1 vccd1 vccd1 _09372_ sky130_fd_sc_hd__a21o_1
X_19552_ clknet_leaf_33_i_clk _00483_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[2\] sky130_fd_sc_hd__dfxtp_1
X_13976_ _06601_ _06600_ _06722_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__a21oi_2
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18503_ rbzero.pov.spi_buffer\[21\] rbzero.pov.spi_buffer\[22\] _02466_ vssd1 vssd1
+ vccd1 vccd1 _02469_ sky130_fd_sc_hd__mux2_1
X_15715_ _06781_ _08267_ _04832_ vssd1 vssd1 vccd1 vccd1 _08398_ sky130_fd_sc_hd__o21a_1
XFILLER_111_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12927_ _05682_ _05683_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__xnor2_1
X_16695_ _09302_ _09303_ vssd1 vssd1 vccd1 vccd1 _09304_ sky130_fd_sc_hd__or2b_1
X_19483_ clknet_leaf_53_i_clk _00429_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-10\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_34_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15646_ _08192_ _08196_ _08194_ vssd1 vssd1 vccd1 vccd1 _08329_ sky130_fd_sc_hd__o21a_1
X_12858_ _05609_ _05467_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__nand2_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18365_ _02422_ vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__clkbuf_1
X_11809_ _03459_ _03469_ net15 vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__mux2_1
X_15577_ _07661_ _08134_ _08260_ _07662_ vssd1 vssd1 vccd1 vccd1 _08261_ sky130_fd_sc_hd__o22ai_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ _05450_ _05545_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__and2_1
XFILLER_14_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ rbzero.wall_tracer.trackDistY\[8\] rbzero.wall_tracer.stepDistY\[8\] vssd1
+ vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__or2_1
XFILLER_187_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14528_ _07196_ _07214_ _07215_ _07200_ vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__a22o_1
XFILLER_175_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18296_ _02381_ vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17247_ _01578_ _01579_ _01580_ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__nand3_1
X_19156__318 clknet_1_1__leaf__02747_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__inv_2
XFILLER_147_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14459_ rbzero.wall_tracer.visualWallDist\[-9\] _06855_ _07144_ rbzero.debug_overlay.playerY\[-9\]
+ _07146_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__a221oi_4
XFILLER_179_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17178_ _03483_ _03458_ _05005_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__and3_1
XFILLER_155_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16129_ _08620_ _08622_ _08619_ vssd1 vssd1 vccd1 vccd1 _08742_ sky130_fd_sc_hd__a21bo_1
XFILLER_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19819_ clknet_leaf_14_i_clk _00750_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_otherx\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_30 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_52 net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_63 net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20525_ clknet_leaf_29_i_clk _01456_ vssd1 vssd1 vccd1 vccd1 gpout4.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_193_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19022__197 clknet_1_1__leaf__02734_ vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__inv_2
X_19096__265 clknet_1_1__leaf__02740_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__inv_2
XFILLER_165_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20456_ net136 _01387_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20387_ net447 _01318_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10140_ rbzero.tex_g0\[62\] rbzero.tex_g0\[61\] _03050_ vssd1 vssd1 vccd1 vccd1 _03128_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10071_ rbzero.tex_g1\[30\] rbzero.tex_g1\[31\] _03084_ vssd1 vssd1 vccd1 vccd1 _03092_
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13830_ _06575_ _06586_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__xor2_1
XFILLER_28_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13761_ _06488_ _06490_ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__xnor2_1
X_10973_ rbzero.tex_r0\[51\] _03696_ _03697_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__and3_1
XFILLER_55_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15500_ _08166_ _08168_ vssd1 vssd1 vccd1 vccd1 _08184_ sky130_fd_sc_hd__nor2_1
XFILLER_44_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12712_ _05468_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__clkbuf_4
X_16480_ _08954_ _09076_ vssd1 vssd1 vccd1 vccd1 _09090_ sky130_fd_sc_hd__nor2_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _06440_ _06443_ _06445_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__and3_1
XFILLER_188_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15431_ _07999_ _08001_ _07998_ vssd1 vssd1 vccd1 vccd1 _08116_ sky130_fd_sc_hd__a21o_1
X_12643_ _05358_ _05361_ _05338_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__mux2_1
XFILLER_54_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18150_ _02291_ vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__clkbuf_2
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15362_ _07940_ _08047_ vssd1 vssd1 vccd1 vccd1 _08048_ sky130_fd_sc_hd__xor2_4
XFILLER_54_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12574_ _05116_ _05240_ _05311_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__mux2_1
X_17101_ _09704_ _09705_ vssd1 vssd1 vccd1 vccd1 _09706_ sky130_fd_sc_hd__and2_1
XFILLER_178_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14313_ _03491_ rbzero.wall_tracer.stepDistY\[-8\] _06906_ vssd1 vssd1 vccd1 vccd1
+ _07001_ sky130_fd_sc_hd__a21oi_1
XFILLER_168_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11525_ _04236_ _04239_ _03764_ _04307_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__a2bb2o_1
X_18081_ _02244_ _02224_ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__or2_2
X_15293_ _07273_ _07092_ vssd1 vssd1 vccd1 vccd1 _07979_ sky130_fd_sc_hd__or2_1
X_17032_ _09007_ _09036_ vssd1 vssd1 vccd1 vccd1 _09637_ sky130_fd_sc_hd__nor2_1
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14244_ _04948_ _06926_ _06930_ _06931_ vssd1 vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__a2bb2o_2
X_11456_ _03540_ _04237_ _04238_ _03997_ _03764_ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__a311o_1
XFILLER_125_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10407_ rbzero.tex_b0\[63\] rbzero.tex_b0\[62\] _03188_ vssd1 vssd1 vccd1 vccd1 _03268_
+ sky130_fd_sc_hd__mux2_1
XFILLER_171_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14175_ _04831_ _06631_ _06862_ vssd1 vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__a21o_1
X_11387_ _04169_ _04170_ _03823_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__mux2_1
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13126_ _05521_ _05878_ _05881_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__o21ai_1
XFILLER_112_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10338_ _03072_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__clkbuf_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _05812_ _05813_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__and2_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ rbzero.pov.spi_buffer\[21\] rbzero.pov.ready_buffer\[21\] _02164_ vssd1 vssd1
+ vccd1 vccd1 _02167_ sky130_fd_sc_hd__mux2_1
X_10269_ rbzero.tex_g0\[1\] rbzero.tex_g0\[0\] _03188_ vssd1 vssd1 vccd1 vccd1 _03196_
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12008_ _04779_ _03913_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__nor2_1
XFILLER_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17865_ _02113_ _02105_ _02122_ _02123_ vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__a31o_1
XFILLER_66_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xnet99_2 clknet_1_0__leaf__04486_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__inv_2
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19604_ clknet_leaf_35_i_clk _00535_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_16816_ _09400_ _09401_ vssd1 vssd1 vccd1 vccd1 _09423_ sky130_fd_sc_hd__or2b_1
XFILLER_93_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17796_ _08458_ _02052_ _02053_ _02061_ vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__a31o_1
XFILLER_4_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19535_ clknet_leaf_66_i_clk _00006_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_16747_ _09258_ _09259_ _09261_ vssd1 vssd1 vccd1 vccd1 _09355_ sky130_fd_sc_hd__a21o_1
XFILLER_34_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13959_ _06601_ _06572_ _06621_ vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__a21oi_1
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16678_ _09284_ _09285_ vssd1 vssd1 vccd1 vccd1 _09287_ sky130_fd_sc_hd__and2_1
X_19466_ clknet_leaf_58_i_clk _00412_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15629_ _08299_ _08302_ _08297_ vssd1 vssd1 vccd1 vccd1 _08312_ sky130_fd_sc_hd__a21bo_1
X_19397_ _08460_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__buf_4
XFILLER_50_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18348_ _02409_ vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18279_ rbzero.spi_registers.spi_buffer\[1\] rbzero.spi_registers.new_floor\[1\]
+ _02370_ vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__mux2_1
X_20310_ net370 _01241_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput50 i_tex_in[3] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__buf_4
XFILLER_162_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20241_ net301 _01172_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20172_ net232 _01103_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09983_ _03045_ vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19210__367 clknet_1_0__leaf__02752_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__inv_2
XFILLER_130_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19104__272 clknet_1_0__leaf__02741_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__inv_2
XFILLER_194_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11310_ rbzero.debug_overlay.facingY\[-4\] _04089_ _04090_ rbzero.debug_overlay.facingY\[-8\]
+ _04094_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__a221o_1
X_20508_ clknet_leaf_30_i_clk _01439_ vssd1 vssd1 vccd1 vccd1 gpout0.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12290_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] rbzero.wall_tracer.rayAddendX\[5\]
+ rbzero.debug_overlay.facingX\[-3\] vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__o211a_1
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11241_ gpout0.vpos\[5\] _03523_ _03524_ _03517_ _04025_ vssd1 vssd1 vccd1 vccd1
+ _04026_ sky130_fd_sc_hd__o221a_1
X_20439_ net499 _01370_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11172_ _03648_ _03943_ _03947_ _03687_ _03956_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__a311o_1
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10123_ _03119_ vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15980_ rbzero.wall_tracer.trackDistX\[-1\] rbzero.wall_tracer.stepDistX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _08594_ sky130_fd_sc_hd__nand2_1
XFILLER_94_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14931_ _06872_ _07119_ _07101_ _07048_ vssd1 vssd1 vccd1 vccd1 _07619_ sky130_fd_sc_hd__or4_1
X_10054_ rbzero.tex_g1\[38\] rbzero.tex_g1\[39\] _03073_ vssd1 vssd1 vccd1 vccd1 _03083_
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14862_ _07539_ _07549_ vssd1 vssd1 vccd1 vccd1 _07550_ sky130_fd_sc_hd__xnor2_1
X_17650_ _01920_ _01925_ _01926_ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16601_ _09208_ _09209_ vssd1 vssd1 vccd1 vccd1 _09210_ sky130_fd_sc_hd__nor2_1
X_13813_ _06284_ _06568_ _06569_ vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__a21o_1
X_17581_ _01785_ rbzero.wall_tracer.rayAddendY\[8\] vssd1 vssd1 vccd1 vccd1 _01867_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_90_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14793_ _07434_ _07437_ vssd1 vssd1 vccd1 vccd1 _07481_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16532_ _08133_ vssd1 vssd1 vccd1 vccd1 _09142_ sky130_fd_sc_hd__buf_2
X_19320_ _02805_ _02806_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__or2_1
X_13744_ _06498_ _06499_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__nand2_1
XFILLER_17_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10956_ rbzero.tex_r0\[39\] rbzero.tex_r0\[38\] _03662_ vssd1 vssd1 vccd1 vccd1 _03742_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16463_ _09071_ _09073_ vssd1 vssd1 vccd1 vccd1 _09074_ sky130_fd_sc_hd__xor2_2
X_13675_ _06427_ _06429_ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__nor2_1
X_10887_ _03606_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__buf_6
XFILLER_43_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15414_ _07973_ _08097_ _08098_ vssd1 vssd1 vccd1 vccd1 _08099_ sky130_fd_sc_hd__o21ai_1
X_18202_ _02319_ _02321_ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__or2_1
X_12626_ _05244_ _05276_ _05297_ _05382_ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__a31o_1
XFILLER_188_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16394_ _08973_ _09004_ vssd1 vssd1 vccd1 vccd1 _09005_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18133_ _03871_ _02263_ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__nand2_1
X_15345_ _08028_ _08030_ vssd1 vssd1 vccd1 vccd1 _08031_ sky130_fd_sc_hd__xnor2_2
X_12557_ _05238_ _05242_ _05313_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__mux2_1
XFILLER_89_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11508_ rbzero.tex_g1\[33\] rbzero.tex_g1\[32\] _03727_ vssd1 vssd1 vccd1 vccd1 _04291_
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18064_ rbzero.spi_registers.spi_buffer\[8\] rbzero.spi_registers.spi_buffer\[7\]
+ _02227_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__mux2_1
X_15276_ _07011_ _07961_ vssd1 vssd1 vccd1 vccd1 _07962_ sky130_fd_sc_hd__nor2_1
XFILLER_117_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12488_ _05215_ _05219_ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__or2_1
X_17015_ _09615_ _09619_ _09620_ vssd1 vssd1 vccd1 vccd1 _09621_ sky130_fd_sc_hd__a21oi_1
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14227_ rbzero.debug_overlay.playerX\[-8\] _06914_ _04838_ vssd1 vssd1 vccd1 vccd1
+ _06915_ sky130_fd_sc_hd__a21oi_1
X_11439_ _03685_ _04214_ _04222_ _03718_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__a31o_1
XFILLER_125_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14158_ net72 rbzero.wall_tracer.wall\[1\] _04827_ vssd1 vssd1 vccd1 vccd1 _06848_
+ sky130_fd_sc_hd__and3_1
XFILLER_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _05479_ _05474_ _05480_ _05609_ vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__o22a_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ rbzero.wall_tracer.visualWallDist\[5\] _03495_ _06785_ rbzero.wall_tracer.trackDistY\[5\]
+ _03497_ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__o221a_1
XFILLER_65_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917_ rbzero.pov.spi_buffer\[13\] rbzero.pov.ready_buffer\[13\] _02153_ vssd1 vssd1
+ vccd1 vccd1 _02158_ sky130_fd_sc_hd__mux2_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18897_ _02257_ _03907_ _02713_ vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__or3_1
XFILLER_117_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17848_ _02107_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[3\]
+ _02108_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__a211o_1
XFILLER_54_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17779_ _02044_ _02045_ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__nor2_1
XFILLER_93_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19518_ clknet_leaf_54_i_clk _00464_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19449_ gpout4.clk_div\[1\] gpout4.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__nand2_1
XFILLER_50_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20224_ net284 _01155_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20155_ net215 _01086_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[2\] sky130_fd_sc_hd__dfxtp_1
X_19134__298 clknet_1_0__leaf__02745_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__inv_2
X_09966_ _03036_ vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20086_ clknet_leaf_84_i_clk _01017_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _03000_ vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _03591_ _03592_ _03595_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__o21bai_2
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ net16 vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__inv_2
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10741_ gpout0.hpos\[1\] vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__buf_2
XFILLER_201_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13460_ _06198_ _06201_ _06216_ vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__nand3_1
X_10672_ _02900_ _03466_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__or2_2
XFILLER_139_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12411_ _03388_ rbzero.wall_tracer.visualWallDist\[9\] _03480_ _03489_ vssd1 vssd1
+ vccd1 vccd1 _05168_ sky130_fd_sc_hd__or4_1
XFILLER_159_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13391_ _05503_ _05992_ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__or2_1
XFILLER_182_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15130_ rbzero.debug_overlay.playerY\[-9\] rbzero.debug_overlay.playerX\[-9\] _06850_
+ vssd1 vssd1 vccd1 vccd1 _07818_ sky130_fd_sc_hd__mux2_1
XFILLER_166_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12342_ _03479_ _04904_ _05098_ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__a21o_1
XFILLER_154_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15061_ _07148_ _07748_ vssd1 vssd1 vccd1 vccd1 _07749_ sky130_fd_sc_hd__or2_1
X_12273_ rbzero.debug_overlay.facingX\[-1\] rbzero.wall_tracer.rayAddendX\[7\] vssd1
+ vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__or2_1
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14012_ _06754_ vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11224_ _03900_ _03901_ _03464_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18820_ _04828_ vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__buf_2
X_11155_ rbzero.tex_r1\[46\] _03620_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__or2_1
XFILLER_95_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10106_ _03110_ vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18751_ rbzero.pov.ready_buffer\[58\] vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__inv_2
X_11086_ rbzero.map_overlay.i_otherx\[3\] vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__inv_2
X_15963_ rbzero.wall_tracer.trackDistX\[-2\] rbzero.wall_tracer.stepDistX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _08579_ sky130_fd_sc_hd__nand2_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17702_ _01972_ rbzero.wall_tracer.rayAddendX\[0\] vssd1 vssd1 vccd1 vccd1 _01974_
+ sky130_fd_sc_hd__and2_1
X_10037_ _03074_ vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__clkbuf_1
X_14914_ _07549_ _07582_ _07580_ vssd1 vssd1 vccd1 vccd1 _07602_ sky130_fd_sc_hd__o21a_1
X_18682_ rbzero.debug_overlay.playerX\[4\] _02570_ _02411_ vssd1 vssd1 vccd1 vccd1
+ _02576_ sky130_fd_sc_hd__o21ai_1
XFILLER_75_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15894_ rbzero.wall_tracer.trackDistX\[-10\] rbzero.wall_tracer.stepDistX\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _08518_ sky130_fd_sc_hd__or2_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17633_ _01911_ vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__clkbuf_1
X_14845_ _07119_ _07005_ vssd1 vssd1 vccd1 vccd1 _07533_ sky130_fd_sc_hd__nor2_1
XFILLER_29_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_5_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17564_ rbzero.wall_tracer.rayAddendY\[6\] _08447_ _01851_ _01714_ vssd1 vssd1 vccd1
+ vccd1 _01852_ sky130_fd_sc_hd__a22o_1
X_14776_ _07433_ _07440_ _07442_ vssd1 vssd1 vccd1 vccd1 _07464_ sky130_fd_sc_hd__and3_1
X_11988_ net39 _04731_ _04724_ net49 vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__a22o_1
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18385__29 clknet_1_0__leaf__02434_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__inv_2
X_19303_ _02791_ _02792_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__xnor2_1
X_16515_ _09123_ _09124_ vssd1 vssd1 vccd1 vccd1 _09125_ sky130_fd_sc_hd__nor2_1
X_13727_ _06103_ _06230_ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__nor2_1
XFILLER_1_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10939_ _03661_ _03722_ _03724_ _03689_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__o211a_1
X_17495_ _01786_ rbzero.wall_tracer.rayAddendY\[2\] vssd1 vssd1 vccd1 vccd1 _01787_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_56_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16446_ _09055_ _09056_ vssd1 vssd1 vccd1 vccd1 _09057_ sky130_fd_sc_hd__nor2_1
X_13658_ _06413_ _06414_ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__nor2_1
XFILLER_108_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _05178_ _05348_ _05324_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__mux2_1
X_19165_ clknet_1_1__leaf__02743_ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__buf_1
X_16377_ _08000_ _07123_ _07333_ _07787_ vssd1 vssd1 vccd1 vccd1 _08988_ sky130_fd_sc_hd__or4_1
XFILLER_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13589_ _05503_ _06156_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__nor2_1
XFILLER_173_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18116_ rbzero.spi_registers.new_other\[7\] _02264_ _02267_ _02266_ vssd1 vssd1 vccd1
+ vccd1 _00751_ sky130_fd_sc_hd__o211a_1
X_15328_ _06771_ _07893_ vssd1 vssd1 vccd1 vccd1 _08014_ sky130_fd_sc_hd__nand2_1
XFILLER_157_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15259_ _07007_ _07332_ _07835_ vssd1 vssd1 vccd1 vccd1 _07945_ sky130_fd_sc_hd__o21bai_1
X_18047_ _02226_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__clkbuf_4
XFILLER_144_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09820_ _02958_ vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19998_ clknet_leaf_93_i_clk _00929_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09751_ _02922_ vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19216__373 clknet_1_1__leaf__02752_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__inv_2
XFILLER_104_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20207_ net267 _01138_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09949_ _03027_ vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__clkbuf_1
X_20138_ clknet_leaf_85_i_clk _01069_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ _05675_ _05676_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20069_ clknet_leaf_67_i_clk _01000_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11911_ _04669_ _04685_ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__and2_1
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _05477_ _05549_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__nand2_2
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _07292_ _07317_ vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__xor2_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ net14 _04617_ net10 net11 vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__and4b_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _07040_ _07247_ _07248_ vssd1 vssd1 vccd1 vccd1 _07249_ sky130_fd_sc_hd__a21bo_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ net8 net7 net62 _04514_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__or4b_1
XFILLER_198_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _07530_ _08018_ _08911_ vssd1 vssd1 vccd1 vccd1 _08912_ sky130_fd_sc_hd__or3b_1
X_13512_ _06255_ _06267_ _06268_ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__a21oi_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ rbzero.wall_tracer.state\[10\] _03510_ _03498_ vssd1 vssd1 vccd1 vccd1 _00014_
+ sky130_fd_sc_hd__o21a_1
X_17280_ rbzero.wall_tracer.trackDistY\[3\] rbzero.wall_tracer.stepDistY\[3\] vssd1
+ vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__nand2_1
XFILLER_14_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _07168_ _07173_ _07174_ _07176_ _07179_ vssd1 vssd1 vccd1 vccd1 _07180_ sky130_fd_sc_hd__a32oi_4
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16231_ _08735_ _08736_ _08739_ vssd1 vssd1 vccd1 vccd1 _08843_ sky130_fd_sc_hd__o21a_1
X_13443_ _06080_ _06081_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__nand2_1
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10655_ rbzero.map_overlay.i_mapdy\[4\] vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__inv_2
XFILLER_139_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16162_ _08647_ _08773_ _08774_ vssd1 vssd1 vccd1 vccd1 _08775_ sky130_fd_sc_hd__a21bo_1
XFILLER_10_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13374_ _06126_ _06130_ _06124_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__o21a_1
XFILLER_155_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10586_ rbzero.wall_tracer.mapX\[9\] rbzero.wall_tracer.mapX\[8\] rbzero.wall_tracer.mapX\[10\]
+ _03381_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__or4_1
XFILLER_186_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15113_ _07329_ _07338_ _07800_ vssd1 vssd1 vccd1 vccd1 _07801_ sky130_fd_sc_hd__a21oi_4
X_12325_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] vssd1
+ vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__xor2_1
XFILLER_182_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16093_ _08705_ _08706_ vssd1 vssd1 vccd1 vccd1 _08707_ sky130_fd_sc_hd__or2_1
XFILLER_177_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19921_ net150 _00852_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[1\] sky130_fd_sc_hd__dfxtp_1
X_15044_ _06968_ _07141_ vssd1 vssd1 vccd1 vccd1 _07732_ sky130_fd_sc_hd__or2_1
XFILLER_177_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12256_ rbzero.wall_tracer.mapY\[8\] _04929_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11207_ rbzero.tex_r1\[17\] _03660_ _03768_ _03670_ vssd1 vssd1 vccd1 vccd1 _03992_
+ sky130_fd_sc_hd__a31o_1
X_19852_ clknet_leaf_25_i_clk _00783_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12187_ _04948_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__buf_4
XFILLER_122_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18803_ rbzero.debug_overlay.facingY\[-2\] _02645_ vssd1 vssd1 vccd1 vccd1 _02662_
+ sky130_fd_sc_hd__and2_1
XFILLER_110_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11138_ rbzero.tex_r1\[50\] _03767_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__or2_1
XFILLER_122_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19783_ clknet_leaf_81_i_clk _00714_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16995_ _09599_ _09600_ vssd1 vssd1 vccd1 vccd1 _09601_ sky130_fd_sc_hd__nand2_1
XFILLER_77_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18734_ rbzero.debug_overlay.playerY\[2\] _02610_ vssd1 vssd1 vccd1 vccd1 _02615_
+ sky130_fd_sc_hd__nand2_1
X_11069_ rbzero.map_overlay.i_mapdy\[3\] rbzero.map_overlay.i_mapdy\[2\] rbzero.map_overlay.i_mapdy\[1\]
+ rbzero.map_overlay.i_mapdy\[0\] vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__or4_1
X_15946_ rbzero.wall_tracer.trackDistX\[-4\] rbzero.wall_tracer.stepDistX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _08564_ sky130_fd_sc_hd__nand2_1
XFILLER_23_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18665_ rbzero.pov.ready_buffer\[68\] _02411_ _02413_ _02562_ _02543_ vssd1 vssd1
+ vccd1 vccd1 _02563_ sky130_fd_sc_hd__o221a_1
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15877_ rbzero.wall_tracer.mapX\[10\] _08502_ vssd1 vssd1 vccd1 vccd1 _08503_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17616_ _08509_ _04935_ _01896_ _01897_ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__a31o_1
XFILLER_64_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14828_ _07458_ _07500_ _07512_ _07513_ _07515_ vssd1 vssd1 vccd1 vccd1 _07516_ sky130_fd_sc_hd__a32oi_2
X_18596_ _02517_ vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17547_ _01834_ _01835_ _01818_ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__o21a_1
XFILLER_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14759_ _07381_ _07390_ vssd1 vssd1 vccd1 vccd1 _07447_ sky130_fd_sc_hd__xnor2_1
XFILLER_177_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17478_ _01771_ vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__clkbuf_1
X_16429_ _07992_ _09039_ vssd1 vssd1 vccd1 vccd1 _09040_ sky130_fd_sc_hd__nor2_1
XFILLER_34_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09803_ _02949_ vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09734_ _02913_ vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10440_ _03285_ vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10371_ _03249_ vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12110_ _04870_ _04871_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__or2_1
X_13090_ _05837_ _05844_ _05846_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__and3_1
XFILLER_117_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12041_ gpout0.vpos\[0\] gpout0.vpos\[1\] _04790_ vssd1 vssd1 vccd1 vccd1 _04814_
+ sky130_fd_sc_hd__mux2_1
XFILLER_133_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15800_ _08448_ vssd1 vssd1 vccd1 vccd1 _08457_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_70_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_65_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16780_ _09386_ _09387_ vssd1 vssd1 vccd1 vccd1 _09388_ sky130_fd_sc_hd__or2_1
XFILLER_120_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13992_ _05373_ _06678_ _06629_ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__a21oi_1
XFILLER_46_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15731_ _08411_ _08412_ vssd1 vssd1 vccd1 vccd1 _08414_ sky130_fd_sc_hd__nand2_1
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ _05689_ _05695_ _05699_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__o21a_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _08343_ _08344_ vssd1 vssd1 vccd1 vccd1 _08345_ sky130_fd_sc_hd__nor2_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12874_ _05519_ _05522_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__or2b_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.wall_tracer.rayAddendY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_85_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ _07295_ _07300_ vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__xnor2_1
X_11825_ _03906_ _04499_ _03909_ gpout0.vpos\[1\] _04559_ _04552_ vssd1 vssd1 vccd1
+ vccd1 _04602_ sky130_fd_sc_hd__mux4_1
X_15593_ _08137_ _08151_ _08150_ vssd1 vssd1 vccd1 vccd1 _08277_ sky130_fd_sc_hd__a21boi_1
X_18381_ clknet_1_0__leaf__04486_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__buf_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14544_ _06940_ _06970_ vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__nor2_1
X_17332_ rbzero.wall_tracer.trackDistY\[10\] rbzero.wall_tracer.stepDistY\[10\] vssd1
+ vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__nand2_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11756_ net44 _04519_ _04513_ _04533_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__a31o_1
XFILLER_183_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10707_ _03495_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__clkbuf_4
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14475_ _06630_ _06752_ vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__nor2_1
X_17263_ _04963_ _01527_ _01594_ vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__a21oi_1
XFILLER_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11687_ _03718_ _04450_ _04467_ _03537_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__a31o_1
XFILLER_146_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16214_ _08702_ _08703_ _08705_ vssd1 vssd1 vccd1 vccd1 _08827_ sky130_fd_sc_hd__a21oi_1
X_13426_ _06162_ _06163_ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__xnor2_1
X_10638_ rbzero.map_overlay.i_othery\[2\] _03345_ vssd1 vssd1 vccd1 vccd1 _03434_
+ sky130_fd_sc_hd__or2_1
X_17194_ _01530_ _01531_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__and2_1
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16145_ _08756_ _08757_ vssd1 vssd1 vccd1 vccd1 _08758_ sky130_fd_sc_hd__nor2_1
XFILLER_155_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13357_ _06096_ _06113_ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__nand2_1
X_10569_ _03363_ _03353_ _03364_ rbzero.debug_overlay.playerX\[4\] vssd1 vssd1 vccd1
+ vccd1 _03365_ sky130_fd_sc_hd__a22o_1
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12308_ _03489_ _05064_ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__nand2_1
X_16076_ _08687_ _08689_ vssd1 vssd1 vccd1 vccd1 _08690_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_23_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_114_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13288_ _05301_ _06008_ _05954_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__or3_1
XFILLER_64_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15027_ _07097_ _07039_ _07273_ _06940_ vssd1 vssd1 vccd1 vccd1 _07715_ sky130_fd_sc_hd__o22ai_1
X_19904_ clknet_leaf_23_i_clk _00835_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12239_ _04956_ rbzero.wall_tracer.trackDistX\[8\] _04957_ rbzero.wall_tracer.trackDistX\[7\]
+ _05000_ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__a221o_1
XFILLER_190_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19835_ clknet_leaf_4_i_clk _00766_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_38_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_110_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19766_ clknet_leaf_85_i_clk _00697_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16978_ _08896_ _09110_ vssd1 vssd1 vccd1 vccd1 _09584_ sky130_fd_sc_hd__nor2_1
XFILLER_49_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput4 i_gpout0_sel[1] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_6
X_18717_ rbzero.debug_overlay.playerY\[-3\] _02588_ _02602_ _02586_ vssd1 vssd1 vccd1
+ vccd1 _01017_ sky130_fd_sc_hd__o211a_1
XFILLER_83_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15929_ _08540_ _08542_ _08541_ vssd1 vssd1 vccd1 vccd1 _08549_ sky130_fd_sc_hd__o21bai_1
X_19697_ clknet_leaf_79_i_clk _00628_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_36_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18648_ _02534_ _02549_ _02550_ _02356_ vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__o211a_1
XFILLER_64_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18441__80 clknet_1_0__leaf__02439_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__inv_2
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18579_ _02508_ vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20472_ net128 _01403_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09717_ gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__buf_2
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19027__202 clknet_1_1__leaf__02734_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__inv_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _03534_ _04389_ _04391_ _04231_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__o211a_1
XFILLER_187_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12590_ _05274_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__clkbuf_4
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11541_ _04198_ _04318_ _04322_ _03721_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__a211o_1
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14260_ rbzero.debug_overlay.playerX\[-5\] _06887_ _04838_ vssd1 vssd1 vccd1 vccd1
+ _06948_ sky130_fd_sc_hd__a21oi_1
XFILLER_156_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ _03671_ _04250_ _04254_ _03721_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__a211o_1
XFILLER_11_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13211_ _05965_ _05967_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__and2_1
XFILLER_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10423_ _03276_ vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14191_ _06877_ _06878_ vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__and2_1
XFILLER_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13142_ _05894_ _05898_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__xor2_1
XFILLER_3_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19073__244 clknet_1_1__leaf__02738_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__inv_2
X_10354_ _03240_ vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13073_ _05792_ _05794_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__and2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17950_ _02142_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__clkbuf_4
XFILLER_3_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10285_ _03204_ vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16901_ _09428_ _09507_ vssd1 vssd1 vccd1 vccd1 _09508_ sky130_fd_sc_hd__xor2_2
X_12024_ net34 _04779_ _03911_ _04796_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__a31o_1
XFILLER_78_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17881_ rbzero.spi_registers.spi_counter\[5\] _02136_ vssd1 vssd1 vccd1 vccd1 _02137_
+ sky130_fd_sc_hd__and2_1
XFILLER_120_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19620_ clknet_leaf_52_i_clk _00551_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16832_ _09437_ _09438_ vssd1 vssd1 vccd1 vccd1 _09439_ sky130_fd_sc_hd__xor2_1
XFILLER_120_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19551_ clknet_leaf_33_i_clk _00482_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16763_ _09361_ _09370_ vssd1 vssd1 vccd1 vccd1 _09371_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13975_ _06588_ _06587_ vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__and2_1
XFILLER_93_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18502_ _02468_ vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15714_ rbzero.wall_tracer.stepDistY\[10\] vssd1 vssd1 vccd1 vccd1 _08397_ sky130_fd_sc_hd__inv_2
X_12926_ _05600_ _05601_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__xor2_1
X_19482_ clknet_leaf_53_i_clk _00428_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
X_16694_ _09204_ _09189_ _09301_ vssd1 vssd1 vccd1 vccd1 _09303_ sky130_fd_sc_hd__a21o_1
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15645_ _08193_ _08327_ vssd1 vssd1 vccd1 vccd1 _08328_ sky130_fd_sc_hd__xnor2_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12857_ _05612_ _05613_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__xor2_1
XFILLER_62_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18364_ _02417_ _02418_ _02421_ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__and3b_1
XFILLER_61_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11808_ net19 _04584_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__nand2_1
XFILLER_159_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15576_ _07897_ vssd1 vssd1 vccd1 vccd1 _08260_ sky130_fd_sc_hd__buf_2
X_12788_ _05495_ _05433_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__nand2_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _01639_ _09520_ rbzero.wall_tracer.trackDistY\[7\] _01523_ vssd1 vssd1 vccd1
+ vccd1 _00578_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14527_ _07195_ _06906_ _03491_ _07107_ vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__or4_1
X_11739_ clknet_leaf_31_i_clk _04516_ _04513_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__and3_2
X_18295_ rbzero.spi_registers.spi_buffer\[1\] rbzero.spi_registers.new_leak\[1\] _02379_
+ vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__mux2_1
XFILLER_187_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17246_ _01572_ _01574_ _01573_ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__o21bai_1
XFILLER_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14458_ _07145_ _04839_ vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__nor2_1
XFILLER_31_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13409_ _06126_ _06130_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__xnor2_1
X_14389_ _06900_ _06970_ vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__nor2_1
X_17177_ _01514_ _01520_ rbzero.wall_tracer.trackDistX\[10\] _08508_ vssd1 vssd1 vccd1
+ vccd1 _00559_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16128_ _08739_ _08740_ vssd1 vssd1 vccd1 vccd1 _08741_ sky130_fd_sc_hd__and2_1
XFILLER_115_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16059_ _07661_ _07662_ _08018_ _08391_ vssd1 vssd1 vccd1 vccd1 _08673_ sky130_fd_sc_hd__or4_1
XFILLER_142_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19818_ clknet_leaf_2_i_clk _00749_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19749_ clknet_leaf_92_i_clk _00680_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_20 rbzero.debug_overlay.facingX\[-4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_31 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_42 net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20524_ clknet_leaf_29_i_clk _01455_ vssd1 vssd1 vccd1 vccd1 gpout4.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_64 net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20455_ net135 _01386_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20386_ net446 _01317_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10070_ _03091_ vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13760_ _06515_ _06516_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__and2_1
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10972_ rbzero.tex_r0\[49\] rbzero.tex_r0\[48\] _03690_ vssd1 vssd1 vccd1 vccd1 _03758_
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12711_ _05392_ _05467_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__or2_1
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13691_ _06418_ _06417_ _06402_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__o21ai_1
XFILLER_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18420__61 clknet_1_1__leaf__02437_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__inv_2
XFILLER_43_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15430_ _08094_ _08114_ vssd1 vssd1 vccd1 vccd1 _08115_ sky130_fd_sc_hd__xnor2_2
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12642_ _05347_ _05394_ _05398_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__a21oi_1
XFILLER_197_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15361_ _08045_ _08046_ vssd1 vssd1 vccd1 vccd1 _08047_ sky130_fd_sc_hd__xor2_4
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12573_ _05329_ _05299_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17100_ _09629_ _09609_ _09703_ vssd1 vssd1 vccd1 vccd1 _09705_ sky130_fd_sc_hd__nand3_1
XFILLER_184_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11524_ _03719_ _04256_ _04273_ _04289_ _04306_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__o32a_1
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14312_ _06955_ _06998_ _06999_ vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__a21bo_1
X_15292_ _07976_ _07977_ vssd1 vssd1 vccd1 vccd1 _07978_ sky130_fd_sc_hd__and2_1
XFILLER_12_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18080_ _02102_ _02103_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__nand2_1
XFILLER_183_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17031_ _09470_ _09533_ _09468_ vssd1 vssd1 vccd1 vccd1 _09636_ sky130_fd_sc_hd__o21a_1
X_14243_ rbzero.debug_overlay.playerX\[-6\] _06914_ _04839_ vssd1 vssd1 vccd1 vccd1
+ _06931_ sky130_fd_sc_hd__a21oi_1
XFILLER_171_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11455_ rbzero.row_render.texu\[2\] _04198_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__nand2_1
XFILLER_183_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10406_ _03267_ vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18938__122 clknet_1_0__leaf__02725_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__inv_2
X_14174_ _06852_ _06861_ _03491_ vssd1 vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__a21o_1
X_11386_ rbzero.tex_g0\[5\] rbzero.tex_g0\[4\] _03615_ vssd1 vssd1 vccd1 vccd1 _04170_
+ sky130_fd_sc_hd__mux2_1
XFILLER_178_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13125_ _05521_ _05878_ _05881_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__or3_1
XFILLER_113_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10337_ _03231_ vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13056_ _05527_ _05610_ _05811_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__o21ai_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ _02166_ vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__clkbuf_1
X_10268_ _03195_ vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12007_ net36 net37 net38 net65 vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__or4_1
XFILLER_87_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17864_ rbzero.spi_registers.spi_counter\[0\] _02102_ _02103_ _02124_ vssd1 vssd1
+ vccd1 vccd1 _00642_ sky130_fd_sc_hd__o211a_1
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10199_ _03159_ vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19603_ clknet_leaf_35_i_clk _00534_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16815_ rbzero.wall_tracer.trackDistX\[6\] _08553_ _09416_ _09422_ vssd1 vssd1 vccd1
+ vccd1 _00555_ sky130_fd_sc_hd__o22a_1
XFILLER_4_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17795_ rbzero.wall_tracer.rayAddendX\[6\] _08447_ _02060_ _01722_ vssd1 vssd1 vccd1
+ vccd1 _02061_ sky130_fd_sc_hd__a22o_1
XFILLER_94_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19534_ clknet_leaf_62_i_clk _00016_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16746_ _09322_ _09353_ vssd1 vssd1 vccd1 vccd1 _09354_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13958_ _05271_ _06604_ _06606_ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__a21o_1
XFILLER_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18984__164 clknet_1_0__leaf__02729_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__inv_2
XFILLER_179_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12909_ _05561_ _05564_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__xor2_1
X_19465_ clknet_leaf_58_i_clk _00411_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16677_ _09284_ _09285_ vssd1 vssd1 vccd1 vccd1 _09286_ sky130_fd_sc_hd__nor2_1
XFILLER_59_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13889_ _06601_ _06614_ _06644_ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__o21bai_1
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15628_ _08182_ _08306_ _08305_ vssd1 vssd1 vccd1 vccd1 _08311_ sky130_fd_sc_hd__a21o_1
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19396_ rbzero.traced_texVinit\[3\] _08463_ _07929_ _01745_ vssd1 vssd1 vccd1 vccd1
+ _01431_ sky130_fd_sc_hd__a22o_1
XFILLER_15_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18347_ rbzero.spi_registers.new_vinf rbzero.spi_registers.spi_buffer\[0\] _02408_
+ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__mux2_1
X_15559_ _08222_ _08242_ vssd1 vssd1 vccd1 vccd1 _08243_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18278_ _02371_ vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__clkbuf_1
Xinput40 i_mode[1] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_8
X_17229_ rbzero.wall_tracer.trackDistY\[-5\] _01523_ _01565_ _08554_ vssd1 vssd1 vccd1
+ vccd1 _00566_ sky130_fd_sc_hd__o22a_1
XFILLER_190_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput51 i_vec_csb vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__buf_8
XFILLER_174_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20240_ net300 _01171_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09982_ rbzero.tex_r0\[9\] rbzero.tex_r0\[8\] _03039_ vssd1 vssd1 vccd1 vccd1 _03045_
+ sky130_fd_sc_hd__mux2_1
XFILLER_192_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20171_ net231 _01102_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__02749_ clknet_0__02749_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02749_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_171_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19139__303 clknet_1_1__leaf__02745_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__inv_2
XFILLER_193_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20507_ clknet_leaf_43_i_clk _01438_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11240_ _03834_ _03466_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__xor2_1
X_20438_ net498 _01369_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11171_ _03949_ _03951_ _03953_ _03955_ _03679_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__o221a_1
X_20369_ net429 _01300_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_122_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10122_ rbzero.tex_g1\[6\] rbzero.tex_g1\[7\] _03117_ vssd1 vssd1 vccd1 vccd1 _03119_
+ sky130_fd_sc_hd__mux2_1
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14930_ _06872_ _07617_ vssd1 vssd1 vccd1 vccd1 _07618_ sky130_fd_sc_hd__nor2_1
X_10053_ _03082_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19185__345 clknet_1_0__leaf__02749_ vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__inv_2
X_14861_ _06872_ _06970_ _07541_ vssd1 vssd1 vccd1 vccd1 _07549_ sky130_fd_sc_hd__nor3_1
XFILLER_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16600_ _09127_ _09205_ _09207_ vssd1 vssd1 vccd1 vccd1 _09209_ sky130_fd_sc_hd__and3_1
X_13812_ _06281_ _06283_ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__nor2_1
X_17580_ _08458_ _01857_ _01858_ _01866_ vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__a31o_1
X_14792_ _07443_ _07468_ vssd1 vssd1 vccd1 vccd1 _07480_ sky130_fd_sc_hd__xnor2_1
XFILLER_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16531_ _09139_ _09140_ vssd1 vssd1 vccd1 vccd1 _09141_ sky130_fd_sc_hd__nand2_1
XFILLER_28_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10955_ rbzero.tex_r0\[37\] rbzero.tex_r0\[36\] _03709_ vssd1 vssd1 vccd1 vccd1 _03741_
+ sky130_fd_sc_hd__mux2_1
X_13743_ _06498_ _06499_ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__or2_1
XFILLER_17_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16462_ _08846_ _08946_ _09072_ vssd1 vssd1 vccd1 vccd1 _09073_ sky130_fd_sc_hd__a21oi_2
X_10886_ _03661_ _03665_ _03668_ _03671_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__o211a_1
XFILLER_177_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13674_ _06426_ _06430_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__and2_1
X_18201_ rbzero.color_sky\[0\] rbzero.spi_registers.new_sky\[0\] _02320_ vssd1 vssd1
+ vccd1 vccd1 _02321_ sky130_fd_sc_hd__mux2_1
X_15413_ _06857_ _06875_ _07097_ _07084_ vssd1 vssd1 vccd1 vccd1 _08098_ sky130_fd_sc_hd__or4_1
X_12625_ _05219_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__inv_2
X_16393_ _09002_ _09003_ vssd1 vssd1 vccd1 vccd1 _09004_ sky130_fd_sc_hd__nand2_1
XFILLER_106_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18132_ rbzero.spi_registers.new_other\[3\] _02264_ _02276_ _02275_ vssd1 vssd1 vccd1
+ vccd1 _00758_ sky130_fd_sc_hd__o211a_1
XFILLER_185_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15344_ _07891_ _07905_ _08029_ vssd1 vssd1 vccd1 vccd1 _08030_ sky130_fd_sc_hd__a21o_1
X_12556_ _05299_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__clkbuf_4
XFILLER_8_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11507_ rbzero.tex_g1\[35\] rbzero.tex_g1\[34\] _03727_ vssd1 vssd1 vccd1 vccd1 _04290_
+ sky130_fd_sc_hd__mux2_1
XFILLER_129_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18063_ _02235_ vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15275_ _07960_ vssd1 vssd1 vccd1 vccd1 _07961_ sky130_fd_sc_hd__clkbuf_4
XFILLER_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12487_ _05234_ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__or2_2
XFILLER_8_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17014_ rbzero.wall_tracer.state\[1\] vssd1 vssd1 vccd1 vccd1 _09620_ sky130_fd_sc_hd__buf_6
X_11438_ _04179_ _04217_ _04221_ _03624_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__a211o_1
X_14226_ _06887_ vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__buf_4
XFILLER_153_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14157_ _06846_ rbzero.mapdxw\[1\] _06842_ vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__mux2_1
X_11369_ _04151_ _04152_ _03666_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__mux2_1
XFILLER_99_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ _05606_ _05607_ _05608_ _05611_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__o2bb2ai_1
X_18965_ clknet_1_1__leaf__02440_ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__buf_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14088_ rbzero.wall_tracer.trackDistX\[4\] _06788_ _06807_ vssd1 vssd1 vccd1 vccd1
+ _00443_ sky130_fd_sc_hd__o21a_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ _05752_ _05753_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__xor2_1
X_17916_ _02157_ vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__clkbuf_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18896_ _03515_ _02714_ _03906_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__a21o_1
XFILLER_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17847_ _02107_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__o21a_1
XFILLER_82_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17778_ _01972_ _04102_ _02042_ _02043_ vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__nor4_1
XFILLER_148_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19517_ clknet_leaf_50_i_clk _00463_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16729_ _07766_ _09229_ vssd1 vssd1 vccd1 vccd1 _09337_ sky130_fd_sc_hd__nor2_1
XFILLER_81_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19448_ gpout4.clk_div\[0\] net61 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__nor2_1
XFILLER_50_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19379_ _02854_ _02855_ _02856_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__a21o_1
XFILLER_10_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20223_ net283 _01154_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20154_ net214 _01085_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[1\] sky130_fd_sc_hd__dfxtp_1
X_09965_ rbzero.tex_r0\[17\] rbzero.tex_r0\[16\] _03028_ vssd1 vssd1 vccd1 vccd1 _03036_
+ sky130_fd_sc_hd__mux2_1
XFILLER_170_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20085_ clknet_leaf_84_i_clk _01016_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
X_09896_ rbzero.tex_r0\[50\] rbzero.tex_r0\[49\] _02995_ vssd1 vssd1 vccd1 vccd1 _03000_
+ sky130_fd_sc_hd__mux2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10740_ gpout0.hpos\[2\] vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__buf_2
XFILLER_159_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10671_ gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__buf_4
XFILLER_186_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ _05159_ _05166_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__nand2_1
XFILLER_199_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13390_ _06145_ _06146_ vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__or2_1
XFILLER_90_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12341_ rbzero.wall_tracer.visualWallDist\[-4\] _05067_ _03487_ vssd1 vssd1 vccd1
+ vccd1 _05098_ sky130_fd_sc_hd__a21o_1
XFILLER_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15060_ _07747_ vssd1 vssd1 vccd1 vccd1 _07748_ sky130_fd_sc_hd__buf_2
X_12272_ rbzero.debug_overlay.facingX\[0\] rbzero.wall_tracer.rayAddendX\[8\] vssd1
+ vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__or2_1
XFILLER_175_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14011_ rbzero.wall_tracer.stepDistY\[3\] _06753_ _06718_ vssd1 vssd1 vccd1 vccd1
+ _06754_ sky130_fd_sc_hd__mux2_1
XFILLER_181_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11223_ gpout0.vpos\[3\] _03523_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__nor2_1
XFILLER_181_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11154_ _03931_ _03933_ _03935_ _03938_ _03648_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__o221a_1
XFILLER_175_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10105_ rbzero.tex_g1\[14\] rbzero.tex_g1\[15\] _03106_ vssd1 vssd1 vccd1 vccd1 _03110_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18750_ _02588_ _02626_ _03360_ vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__a21o_1
XFILLER_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11085_ rbzero.map_overlay.i_othery\[4\] vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__inv_2
X_15962_ rbzero.wall_tracer.trackDistX\[-2\] rbzero.wall_tracer.stepDistX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _08578_ sky130_fd_sc_hd__or2_1
X_17701_ _01972_ rbzero.wall_tracer.rayAddendX\[0\] vssd1 vssd1 vccd1 vccd1 _01973_
+ sky130_fd_sc_hd__nor2_1
XFILLER_88_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10036_ rbzero.tex_g1\[47\] rbzero.tex_g1\[48\] _03073_ vssd1 vssd1 vccd1 vccd1 _03074_
+ sky130_fd_sc_hd__mux2_1
X_14913_ _07599_ _07600_ vssd1 vssd1 vccd1 vccd1 _07601_ sky130_fd_sc_hd__nor2_1
X_18681_ _02543_ _02574_ _03350_ vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__a21oi_1
X_15893_ _07693_ _07695_ _08516_ vssd1 vssd1 vccd1 vccd1 _08517_ sky130_fd_sc_hd__o21a_1
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17632_ _01910_ rbzero.map_rom.i_row\[4\] _05009_ vssd1 vssd1 vccd1 vccd1 _01911_
+ sky130_fd_sc_hd__mux2_1
X_14844_ _07101_ _06978_ vssd1 vssd1 vccd1 vccd1 _07532_ sky130_fd_sc_hd__nor2_1
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17563_ _01849_ _01850_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__xnor2_1
X_14775_ _07445_ _07462_ vssd1 vssd1 vccd1 vccd1 _07463_ sky130_fd_sc_hd__xor2_1
X_11987_ net69 _04731_ _04724_ _03910_ _04760_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__a221o_1
XFILLER_186_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19302_ _02785_ _02788_ _02786_ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__o21bai_1
X_16514_ _09121_ _09122_ vssd1 vssd1 vccd1 vccd1 _09124_ sky130_fd_sc_hd__and2_1
XFILLER_44_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13726_ _06481_ _06482_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__nand2_1
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10938_ _03677_ _03723_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__or2_1
XFILLER_31_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17494_ _01785_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__clkbuf_4
XFILLER_189_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16445_ _09053_ _09054_ vssd1 vssd1 vccd1 vccd1 _09056_ sky130_fd_sc_hd__and2_1
XFILLER_149_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10869_ rbzero.tex_r0\[3\] rbzero.tex_r0\[2\] _03616_ vssd1 vssd1 vccd1 vccd1 _03655_
+ sky130_fd_sc_hd__mux2_1
XFILLER_176_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13657_ _06370_ _06407_ _06412_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__a21oi_1
XFILLER_158_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12608_ _05158_ _05223_ _05313_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__mux2_1
X_16376_ _08000_ _07333_ vssd1 vssd1 vccd1 vccd1 _08987_ sky130_fd_sc_hd__or2_1
XFILLER_157_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13588_ _06008_ _06230_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__or2_1
XFILLER_158_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18115_ _03430_ _02263_ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__nand2_1
XFILLER_200_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15327_ _06771_ _07893_ vssd1 vssd1 vccd1 vccd1 _08013_ sky130_fd_sc_hd__or2_1
XFILLER_117_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12539_ _05224_ _05226_ _05232_ _05295_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__or4b_1
XFILLER_184_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18046_ _02225_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__buf_2
XFILLER_117_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15258_ _07007_ _07049_ _07332_ _07786_ vssd1 vssd1 vccd1 vccd1 _07944_ sky130_fd_sc_hd__or4_1
XFILLER_32_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14209_ _06852_ _06896_ _03490_ vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__a21oi_1
XFILLER_141_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15189_ _07093_ _07733_ _07736_ _07875_ vssd1 vssd1 vccd1 vccd1 _07876_ sky130_fd_sc_hd__a22o_1
XFILLER_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19997_ clknet_leaf_94_i_clk _00928_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09750_ rbzero.tex_r1\[53\] rbzero.tex_r1\[54\] _02921_ vssd1 vssd1 vccd1 vccd1 _02922_
+ sky130_fd_sc_hd__mux2_1
XFILLER_100_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18879_ _04827_ _02702_ _08439_ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__a21o_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18908__95 clknet_1_0__leaf__02441_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__inv_2
XFILLER_195_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20206_ net266 _01137_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20137_ clknet_leaf_85_i_clk _01068_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_09948_ rbzero.tex_r0\[25\] rbzero.tex_r0\[24\] _03017_ vssd1 vssd1 vccd1 vccd1 _03027_
+ sky130_fd_sc_hd__mux2_1
XFILLER_131_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20068_ clknet_leaf_67_i_clk _00999_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-6\]
+ sky130_fd_sc_hd__dfxtp_2
X_09879_ rbzero.tex_r0\[58\] rbzero.tex_r0\[57\] _02984_ vssd1 vssd1 vccd1 vccd1 _02991_
+ sky130_fd_sc_hd__mux2_1
XFILLER_100_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ net24 net23 vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__nor2_2
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _05506_ _05509_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _04612_ net65 _04615_ _04616_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__a211o_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14560_ _07235_ _07037_ _07025_ vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__or3_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ net8 _04527_ _04539_ _04549_ _04533_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__a311o_1
XFILLER_41_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _06257_ _06266_ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__nor2_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _03506_ rbzero.wall_tracer.state\[14\] vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__and2b_1
XFILLER_199_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ _07158_ _07167_ _07178_ vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__or3_2
XFILLER_158_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _08762_ _08728_ vssd1 vssd1 vccd1 vccd1 _08842_ sky130_fd_sc_hd__or2b_1
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13442_ _06080_ _06081_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__nor2_1
X_10654_ rbzero.map_overlay.i_mapdy\[1\] _03374_ _03359_ rbzero.map_overlay.i_mapdy\[4\]
+ _03449_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__o221a_1
XFILLER_13_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16161_ _08229_ _07748_ _08366_ vssd1 vssd1 vccd1 vccd1 _08774_ sky130_fd_sc_hd__or3_1
XFILLER_142_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13373_ _06123_ _06129_ _06097_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__a21oi_1
XFILLER_182_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10585_ rbzero.wall_tracer.mapY\[6\] rbzero.wall_tracer.mapY\[9\] rbzero.wall_tracer.mapY\[8\]
+ rbzero.wall_tracer.mapY\[10\] vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__or4_1
XFILLER_103_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15112_ _07291_ _07328_ vssd1 vssd1 vccd1 vccd1 _07800_ sky130_fd_sc_hd__nor2_1
XFILLER_86_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12324_ _03489_ _05078_ _05079_ _05080_ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__o31ai_4
XFILLER_186_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16092_ _08603_ _08704_ vssd1 vssd1 vccd1 vccd1 _08706_ sky130_fd_sc_hd__nor2_1
XFILLER_115_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19920_ net149 _00851_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[0\] sky130_fd_sc_hd__dfxtp_1
X_15043_ _07729_ _07730_ _07139_ _07142_ vssd1 vssd1 vccd1 vccd1 _07731_ sky130_fd_sc_hd__a22o_1
X_12255_ rbzero.map_rom.i_row\[4\] rbzero.wall_tracer.mapY\[5\] rbzero.wall_tracer.mapY\[7\]
+ rbzero.wall_tracer.mapY\[6\] _04923_ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__o41a_1
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11206_ rbzero.tex_r1\[19\] _03664_ _03990_ _03677_ vssd1 vssd1 vccd1 vccd1 _03991_
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19851_ clknet_leaf_24_i_clk _00782_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12186_ _04947_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__buf_4
X_11137_ rbzero.tex_r1\[52\] _03920_ _03618_ _03921_ vssd1 vssd1 vccd1 vccd1 _03922_
+ sky130_fd_sc_hd__a31o_1
XFILLER_123_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18802_ rbzero.pov.ready_buffer\[28\] _02636_ _02661_ _02643_ vssd1 vssd1 vccd1 vccd1
+ _01043_ sky130_fd_sc_hd__o211a_1
X_19782_ clknet_leaf_83_i_clk _00713_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_110_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16994_ _09563_ _09598_ vssd1 vssd1 vccd1 vccd1 _09600_ sky130_fd_sc_hd__or2_1
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18733_ rbzero.debug_overlay.playerY\[2\] _02610_ vssd1 vssd1 vccd1 vccd1 _02614_
+ sky130_fd_sc_hd__or2_1
XFILLER_114_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11068_ gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__inv_2
XFILLER_49_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15945_ rbzero.wall_tracer.trackDistX\[-4\] rbzero.wall_tracer.stepDistX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _08563_ sky130_fd_sc_hd__or2_1
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10019_ _03064_ vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18664_ _02560_ _02561_ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__nand2_1
XFILLER_64_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15876_ rbzero.wall_tracer.mapX\[9\] _07826_ _08501_ vssd1 vssd1 vccd1 vccd1 _08502_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_92_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17615_ _03357_ _09620_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__nor2_1
XFILLER_184_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14827_ _07514_ _07512_ vssd1 vssd1 vccd1 vccd1 _07515_ sky130_fd_sc_hd__xnor2_1
X_18595_ rbzero.pov.spi_buffer\[65\] rbzero.pov.spi_buffer\[66\] _02510_ vssd1 vssd1
+ vccd1 vccd1 _02517_ sky130_fd_sc_hd__mux2_1
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17546_ _01784_ rbzero.debug_overlay.vplaneY\[-3\] vssd1 vssd1 vccd1 vccd1 _01835_
+ sky130_fd_sc_hd__and2_1
X_14758_ _07438_ _07439_ vssd1 vssd1 vccd1 vccd1 _07446_ sky130_fd_sc_hd__xnor2_1
XFILLER_17_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13709_ _06447_ _06448_ _06465_ vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__a21o_1
XFILLER_189_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17477_ rbzero.wall_tracer.rayAddendY\[0\] _01770_ _03509_ vssd1 vssd1 vccd1 vccd1
+ _01771_ sky130_fd_sc_hd__mux2_1
X_14689_ _06932_ _06969_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__nor2_1
XFILLER_20_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16428_ _08260_ vssd1 vssd1 vccd1 vccd1 _09039_ sky130_fd_sc_hd__clkbuf_4
XFILLER_34_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16359_ _08879_ _08968_ _08969_ vssd1 vssd1 vccd1 vccd1 _08970_ sky130_fd_sc_hd__a21oi_1
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18029_ _02216_ vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09802_ rbzero.tex_r1\[28\] rbzero.tex_r1\[29\] _02943_ vssd1 vssd1 vccd1 vccd1 _02949_
+ sky130_fd_sc_hd__mux2_1
XFILLER_119_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09733_ rbzero.tex_r1\[61\] rbzero.tex_r1\[62\] _02910_ vssd1 vssd1 vccd1 vccd1 _02913_
+ sky130_fd_sc_hd__mux2_1
X_19243__17 clknet_1_0__leaf__02755_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__inv_2
XFILLER_28_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10370_ rbzero.tex_b1\[16\] rbzero.tex_b1\[17\] _03243_ vssd1 vssd1 vccd1 vccd1 _03249_
+ sky130_fd_sc_hd__mux2_1
XFILLER_164_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_4_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_152_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12040_ _04792_ _04811_ _04812_ _04808_ net36 vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__a221o_1
XFILLER_137_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18427__67 clknet_1_1__leaf__02438_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__inv_2
XFILLER_120_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13991_ _06690_ _06708_ _06723_ _06735_ _06664_ _06675_ vssd1 vssd1 vccd1 vccd1 _06736_
+ sky130_fd_sc_hd__mux4_2
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15730_ _08411_ _08412_ vssd1 vssd1 vccd1 vccd1 _08413_ sky130_fd_sc_hd__nor2_1
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _05661_ _05698_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__and2_1
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15661_ _08337_ _08338_ _08342_ vssd1 vssd1 vccd1 vccd1 _08344_ sky130_fd_sc_hd__and3_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _05628_ _05629_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__nand2_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17400_ _01699_ vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__clkbuf_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _07141_ _07157_ _07215_ _07299_ vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__o31a_1
X_18380_ _02432_ vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__clkbuf_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _04579_ _04597_ _04600_ _04571_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__o31a_2
X_15592_ _08264_ _08275_ vssd1 vssd1 vccd1 vccd1 _08276_ sky130_fd_sc_hd__xnor2_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ rbzero.wall_tracer.trackDistY\[10\] rbzero.wall_tracer.stepDistY\[10\] vssd1
+ vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__or2_1
XFILLER_121_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _07229_ _07230_ vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__nor2_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _04532_ _04522_ _04515_ _04525_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__and4_1
XFILLER_57_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17262_ _04946_ _01592_ _01593_ _08717_ _01522_ vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__o311a_1
X_10706_ _03494_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__buf_2
XFILLER_187_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14474_ _07161_ vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__inv_2
XFILLER_201_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11686_ _04458_ _04466_ _03687_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__a21o_1
XFILLER_186_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16213_ _08727_ _08825_ vssd1 vssd1 vccd1 vccd1 _08826_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13425_ _06176_ _06180_ _06181_ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__a21o_1
XFILLER_201_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10637_ rbzero.map_overlay.i_othery\[2\] _03345_ vssd1 vssd1 vccd1 vccd1 _03433_
+ sky130_fd_sc_hd__nand2_1
X_17193_ _08509_ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__clkbuf_4
XFILLER_155_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16144_ _08754_ _08755_ vssd1 vssd1 vccd1 vccd1 _08757_ sky130_fd_sc_hd__and2_1
XFILLER_155_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13356_ _06102_ _06112_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__xor2_1
X_10568_ rbzero.map_rom.i_col\[4\] vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__clkinv_2
XFILLER_127_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12307_ _05060_ _05063_ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__xor2_2
X_16075_ _08395_ _08406_ _08688_ vssd1 vssd1 vccd1 vccd1 _08689_ sky130_fd_sc_hd__a21boi_1
XFILLER_115_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10499_ _03316_ vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13287_ _05964_ _06042_ _06043_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__o21a_1
XFILLER_108_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15026_ _06940_ _07039_ _07713_ vssd1 vssd1 vccd1 vccd1 _07714_ sky130_fd_sc_hd__or3_1
X_19903_ clknet_leaf_21_i_clk _00834_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12238_ _04957_ rbzero.wall_tracer.trackDistX\[7\] _04958_ rbzero.wall_tracer.trackDistX\[6\]
+ _04999_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__o221a_1
XFILLER_123_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19050__223 clknet_1_1__leaf__02736_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__inv_2
X_19834_ clknet_leaf_4_i_clk _00765_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12169_ rbzero.wall_tracer.mapY\[5\] _04929_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16977_ _09581_ _09582_ vssd1 vssd1 vccd1 vccd1 _09583_ sky130_fd_sc_hd__nand2_1
X_19765_ clknet_leaf_86_i_clk _00696_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput5 i_gpout0_sel[2] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_4
X_18716_ rbzero.pov.ready_buffer\[50\] _02413_ _02582_ _02601_ vssd1 vssd1 vccd1 vccd1
+ _02602_ sky130_fd_sc_hd__a211o_1
X_15928_ rbzero.wall_tracer.trackDistX\[-6\] rbzero.wall_tracer.stepDistX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _08548_ sky130_fd_sc_hd__nand2_1
X_19696_ clknet_leaf_79_i_clk _00627_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_76_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18647_ rbzero.debug_overlay.playerX\[-5\] _02542_ vssd1 vssd1 vccd1 vccd1 _02550_
+ sky130_fd_sc_hd__or2_1
XFILLER_65_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15859_ _08487_ vssd1 vssd1 vccd1 vccd1 _08489_ sky130_fd_sc_hd__buf_4
XFILLER_92_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18578_ rbzero.pov.spi_buffer\[57\] rbzero.pov.spi_buffer\[58\] _02499_ vssd1 vssd1
+ vccd1 vccd1 _02508_ sky130_fd_sc_hd__mux2_1
XFILLER_51_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17529_ _01757_ rbzero.debug_overlay.vplaneY\[-4\] vssd1 vssd1 vccd1 vccd1 _01819_
+ sky130_fd_sc_hd__nand2_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20471_ net127 _01402_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11540_ _04319_ _04320_ _04321_ _04192_ _04179_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__o221a_1
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11471_ _04251_ _04252_ _04253_ _03917_ _03674_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__o221a_1
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10422_ rbzero.tex_b0\[56\] rbzero.tex_b0\[55\] _03269_ vssd1 vssd1 vccd1 vccd1 _03276_
+ sky130_fd_sc_hd__mux2_1
X_13210_ _05880_ _05928_ _05964_ _05966_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__o22ai_1
X_14190_ rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerY\[-9\] rbzero.debug_overlay.playerY\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _06878_ sky130_fd_sc_hd__o21ai_1
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10353_ rbzero.tex_b1\[24\] rbzero.tex_b1\[25\] _03232_ vssd1 vssd1 vccd1 vccd1 _03240_
+ sky130_fd_sc_hd__mux2_1
X_13141_ _05896_ _05897_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__and2_1
XFILLER_87_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13072_ _05827_ _05828_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__nor2_1
X_10284_ rbzero.tex_b1\[57\] rbzero.tex_b1\[58\] _03199_ vssd1 vssd1 vccd1 vccd1 _03204_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16900_ _09505_ _09506_ vssd1 vssd1 vccd1 vccd1 _09507_ sky130_fd_sc_hd__nand2_1
X_12023_ net42 _04791_ _04793_ _04795_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__a211o_1
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17880_ _02123_ _02133_ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__nor2_1
X_16831_ _09324_ _09327_ _09326_ vssd1 vssd1 vccd1 vccd1 _09438_ sky130_fd_sc_hd__a21boi_1
XFILLER_120_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19550_ clknet_leaf_32_i_clk _00481_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[0\] sky130_fd_sc_hd__dfxtp_2
X_16762_ _09368_ _09369_ vssd1 vssd1 vccd1 vccd1 _09370_ sky130_fd_sc_hd__nor2_1
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13974_ _06676_ vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__inv_2
XFILLER_93_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18501_ rbzero.pov.spi_buffer\[20\] rbzero.pov.spi_buffer\[21\] _02466_ vssd1 vssd1
+ vccd1 vccd1 _02468_ sky130_fd_sc_hd__mux2_1
X_15713_ _04841_ rbzero.wall_tracer.stepDistX\[10\] vssd1 vssd1 vccd1 vccd1 _08396_
+ sky130_fd_sc_hd__nor2_1
XFILLER_19_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12925_ _05680_ _05664_ _05681_ _05679_ _05678_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__o32a_1
X_19481_ clknet_leaf_50_i_clk _00427_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_16693_ _09204_ _09189_ _09301_ vssd1 vssd1 vccd1 vccd1 _09302_ sky130_fd_sc_hd__and3_1
XFILLER_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15644_ _08209_ _08325_ _08326_ vssd1 vssd1 vccd1 vccd1 _08327_ sky130_fd_sc_hd__a21oi_1
XFILLER_46_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _05536_ _05582_ _05537_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__o21ai_1
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _02414_ _02420_ _02415_ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__a21boi_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ net16 net17 net18 vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__a21o_1
X_15575_ _07617_ _07646_ _07757_ _07897_ vssd1 vssd1 vccd1 vccd1 _08259_ sky130_fd_sc_hd__or4_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _05540_ _05543_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__xnor2_2
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _08512_ _01638_ _01527_ vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__a21oi_1
XFILLER_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _06906_ _07107_ _06985_ _06787_ vssd1 vssd1 vccd1 vccd1 _07214_ sky130_fd_sc_hd__and4bb_1
XFILLER_186_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11738_ net3 net4 vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__and2b_1
X_18294_ _02380_ vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17245_ rbzero.wall_tracer.trackDistY\[-2\] rbzero.wall_tracer.stepDistY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__nand2_1
XFILLER_175_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14457_ rbzero.debug_overlay.playerX\[-9\] vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__clkinv_2
XFILLER_70_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11669_ _04441_ _04449_ _03685_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__a21o_1
XFILLER_30_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13408_ _06142_ _06154_ _06164_ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__o21ai_1
X_17176_ _08524_ _01518_ _01519_ _08507_ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__o31a_1
XFILLER_190_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14388_ _06876_ _07075_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__nor2_2
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16127_ _08737_ _08738_ vssd1 vssd1 vccd1 vccd1 _08740_ sky130_fd_sc_hd__or2_1
X_13339_ _05997_ _06095_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__xor2_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16058_ _07877_ _08260_ vssd1 vssd1 vccd1 vccd1 _08672_ sky130_fd_sc_hd__nor2_1
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18915__101 clknet_1_0__leaf__02723_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__inv_2
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15009_ _07525_ _07573_ vssd1 vssd1 vccd1 vccd1 _07697_ sky130_fd_sc_hd__nor2_1
XFILLER_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19817_ clknet_leaf_2_i_clk _00748_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18406__48 clknet_1_0__leaf__02436_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__inv_2
X_19748_ clknet_leaf_92_i_clk _00679_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19679_ clknet_leaf_80_i_clk _00610_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18961__143 clknet_1_1__leaf__02727_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__inv_2
XFILLER_127_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_10 _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 rbzero.debug_overlay.playerY\[-9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_32 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_43 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20523_ clknet_leaf_41_i_clk _01454_ vssd1 vssd1 vccd1 vccd1 gpout3.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_54 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_65 net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20454_ net134 _01385_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19057__229 clknet_1_1__leaf__02737_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__inv_2
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20385_ net445 _01316_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_84_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_133_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10971_ _03755_ _03756_ _03693_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__mux2_1
XFILLER_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12710_ _05466_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__buf_4
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13690_ _06418_ _06402_ _06417_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_22_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12641_ _05395_ _05396_ _05397_ _05333_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__a211o_1
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15360_ _07796_ _07923_ _07921_ vssd1 vssd1 vccd1 vccd1 _08046_ sky130_fd_sc_hd__a21oi_2
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12572_ _05285_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__clkbuf_4
XFILLER_196_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14311_ _06949_ _06954_ _06966_ _06977_ vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__or4_1
X_11523_ _03685_ _04297_ _04305_ _03718_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__a31o_1
XFILLER_141_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15291_ _07972_ _07270_ _07975_ vssd1 vssd1 vccd1 vccd1 _07977_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_37_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17030_ _09545_ _09556_ _09555_ vssd1 vssd1 vccd1 vccd1 _09635_ sky130_fd_sc_hd__a21o_1
XFILLER_156_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14242_ _06914_ _06929_ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__or2_1
XFILLER_156_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11454_ rbzero.row_render.texu\[2\] _04198_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__or2_1
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10405_ net49 rbzero.tex_b0\[63\] _03188_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__mux2_1
X_11385_ rbzero.tex_g0\[7\] rbzero.tex_g0\[6\] _03615_ vssd1 vssd1 vccd1 vccd1 _04169_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14173_ rbzero.wall_tracer.rayAddendY\[-3\] rbzero.wall_tracer.rayAddendX\[-3\] _06849_
+ vssd1 vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__mux2_1
XFILLER_178_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13124_ _05878_ _05880_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__xnor2_1
XFILLER_194_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10336_ rbzero.tex_b1\[32\] rbzero.tex_b1\[33\] _03221_ vssd1 vssd1 vccd1 vccd1 _03231_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10267_ rbzero.tex_g0\[2\] rbzero.tex_g0\[1\] _03188_ vssd1 vssd1 vccd1 vccd1 _03195_
+ sky130_fd_sc_hd__mux2_1
X_13055_ _05527_ _05610_ _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__or3_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17932_ rbzero.pov.spi_buffer\[20\] rbzero.pov.ready_buffer\[20\] _02164_ vssd1 vssd1
+ vccd1 vccd1 _02166_ sky130_fd_sc_hd__mux2_1
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12006_ net33 vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__buf_2
XFILLER_121_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17863_ _02104_ _02122_ _02123_ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__a21o_1
X_10198_ rbzero.tex_g0\[35\] rbzero.tex_g0\[34\] _03155_ vssd1 vssd1 vccd1 vccd1 _03159_
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19602_ clknet_leaf_35_i_clk _00533_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16814_ _08562_ _09420_ _09421_ _08487_ vssd1 vssd1 vccd1 vccd1 _09422_ sky130_fd_sc_hd__a31o_1
X_17794_ _02058_ _02059_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16745_ _09351_ _09352_ vssd1 vssd1 vccd1 vccd1 _09353_ sky130_fd_sc_hd__nand2_1
X_19533_ clknet_leaf_66_i_clk _00005_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13957_ _06706_ vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__clkbuf_1
X_19162__324 clknet_1_1__leaf__02747_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__inv_2
X_12908_ _05567_ _05568_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__xnor2_1
X_19464_ clknet_leaf_57_i_clk _00410_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16676_ _09164_ _09171_ _09169_ vssd1 vssd1 vccd1 vccd1 _09285_ sky130_fd_sc_hd__a21oi_2
XFILLER_146_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13888_ _05324_ _06611_ vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__nor2_1
XFILLER_179_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18415_ clknet_1_1__leaf__02433_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__buf_1
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15627_ rbzero.wall_tracer.texu\[4\] _06853_ _08309_ _08310_ _03498_ vssd1 vssd1
+ vccd1 vccd1 _00479_ sky130_fd_sc_hd__o221a_1
X_12839_ _05590_ _05595_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__xnor2_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19395_ rbzero.traced_texVinit\[2\] _08463_ _07808_ _01745_ vssd1 vssd1 vccd1 vccd1
+ _01430_ sky130_fd_sc_hd__a22o_1
XFILLER_146_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18346_ _02107_ _01658_ _02907_ _02399_ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__and4_1
X_15558_ _08240_ _08241_ vssd1 vssd1 vccd1 vccd1 _08242_ sky130_fd_sc_hd__nand2_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14509_ _07194_ _07196_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__nor2_1
X_18277_ rbzero.spi_registers.spi_buffer\[0\] rbzero.spi_registers.new_floor\[0\]
+ _02370_ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__mux2_1
X_15489_ _08063_ _08173_ vssd1 vssd1 vccd1 vccd1 _08174_ sky130_fd_sc_hd__xor2_4
XFILLER_147_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17228_ _01534_ _01563_ _01564_ _01526_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__a31o_1
Xinput30 i_gpout4_sel[3] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_4
Xinput41 i_mode[2] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_4
Xinput52 i_vec_mosi vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_4
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17159_ _01498_ _01502_ vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__xnor2_1
X_20170_ net230 _01101_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[17\] sky130_fd_sc_hd__dfxtp_1
X_09981_ _03044_ vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__02748_ clknet_0__02748_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02748_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_157_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20506_ clknet_leaf_42_i_clk _01437_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20437_ net497 _01368_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11170_ rbzero.tex_r1\[32\] _03660_ _03733_ _03954_ vssd1 vssd1 vccd1 vccd1 _03955_
+ sky130_fd_sc_hd__a31o_1
X_20368_ net428 _01299_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10121_ _03118_ vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20299_ net359 _01230_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10052_ rbzero.tex_g1\[39\] rbzero.tex_g1\[40\] _03073_ vssd1 vssd1 vccd1 vccd1 _03082_
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19111__278 clknet_1_0__leaf__02742_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__inv_2
XFILLER_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14860_ _07513_ _07515_ vssd1 vssd1 vccd1 vccd1 _07548_ sky130_fd_sc_hd__xnor2_1
XFILLER_57_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13811_ _06333_ _06566_ _06567_ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__a21o_1
X_18968__149 clknet_1_1__leaf__02728_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__inv_2
XFILLER_35_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14791_ _07427_ _07470_ vssd1 vssd1 vccd1 vccd1 _07479_ sky130_fd_sc_hd__xor2_2
XFILLER_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16530_ _09016_ _08134_ _09039_ _09014_ vssd1 vssd1 vccd1 vccd1 _09140_ sky130_fd_sc_hd__o22ai_1
XFILLER_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13742_ _06103_ _06230_ _06483_ _06481_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__o31a_1
XFILLER_17_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10954_ _03739_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__buf_6
XFILLER_71_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16461_ _08943_ _08945_ vssd1 vssd1 vccd1 vccd1 _09072_ sky130_fd_sc_hd__nor2_1
XFILLER_71_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13673_ _06427_ _06429_ vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__xor2_1
X_10885_ _03670_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__buf_4
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18200_ rbzero.spi_registers.got_new_sky _02261_ vssd1 vssd1 vccd1 vccd1 _02320_
+ sky130_fd_sc_hd__and2_2
X_15412_ _06858_ _07097_ vssd1 vssd1 vccd1 vccd1 _08097_ sky130_fd_sc_hd__nor2_1
XFILLER_176_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12624_ _05377_ _05379_ _05380_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__mux2_1
X_16392_ _08905_ _08974_ _09001_ vssd1 vssd1 vccd1 vccd1 _09003_ sky130_fd_sc_hd__nand3_1
X_18131_ _03873_ _02263_ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__nand2_1
X_15343_ _07904_ _07903_ vssd1 vssd1 vccd1 vccd1 _08029_ sky130_fd_sc_hd__and2b_1
XFILLER_19_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12555_ _05212_ _05217_ _05311_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__mux2_1
X_19005__183 clknet_1_0__leaf__02731_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__inv_2
XFILLER_185_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11506_ _03648_ _04280_ _04284_ _04288_ _03688_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__o221a_1
XFILLER_145_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18062_ rbzero.spi_registers.spi_buffer\[7\] rbzero.spi_registers.spi_buffer\[6\]
+ _02227_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__mux2_1
XFILLER_106_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15274_ _07959_ vssd1 vssd1 vccd1 vccd1 _07960_ sky130_fd_sc_hd__buf_2
XFILLER_157_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12486_ _05238_ _05240_ _05242_ _05116_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__or4b_2
XFILLER_89_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17013_ _09408_ _09409_ _09616_ _09517_ _09618_ vssd1 vssd1 vccd1 vccd1 _09619_ sky130_fd_sc_hd__a41o_2
X_14225_ _06887_ _06912_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__or2_1
XFILLER_171_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11437_ _03656_ _04218_ _04219_ _04220_ _03606_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__o221a_1
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14156_ rbzero.mapdyw\[1\] _06839_ _06840_ _03419_ vssd1 vssd1 vccd1 vccd1 _06846_
+ sky130_fd_sc_hd__a22o_1
XFILLER_99_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11368_ rbzero.tex_g0\[23\] rbzero.tex_g0\[22\] _03709_ vssd1 vssd1 vccd1 vccd1 _04152_
+ sky130_fd_sc_hd__mux2_1
XFILLER_180_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13107_ _05606_ _05861_ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__a21o_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _03222_ vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__clkbuf_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ rbzero.wall_tracer.visualWallDist\[4\] _06796_ _06785_ rbzero.wall_tracer.trackDistY\[4\]
+ _06797_ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__o221a_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11299_ _04067_ _04082_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__nor2_4
XFILLER_79_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13038_ _05792_ _05794_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__nor2_1
X_17915_ rbzero.pov.spi_buffer\[12\] rbzero.pov.ready_buffer\[12\] _02153_ vssd1 vssd1
+ vccd1 vccd1 _02157_ sky130_fd_sc_hd__mux2_1
XFILLER_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18895_ _03907_ _02713_ _02717_ vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__o21a_1
XFILLER_117_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17846_ rbzero.spi_registers.spi_cmd\[0\] vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__clkbuf_2
XFILLER_93_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14989_ _07668_ _07671_ _07674_ vssd1 vssd1 vccd1 vccd1 _07677_ sky130_fd_sc_hd__or3_1
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17777_ _01972_ _04102_ _02042_ _02043_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__o22a_1
XFILLER_187_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19516_ clknet_leaf_50_i_clk _00462_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16728_ _08896_ _08889_ _09250_ _09248_ vssd1 vssd1 vccd1 vccd1 _09336_ sky130_fd_sc_hd__o31a_1
XFILLER_35_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16659_ _09158_ _09159_ _09156_ vssd1 vssd1 vccd1 vccd1 _09268_ sky130_fd_sc_hd__a21o_1
X_19447_ _02895_ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19378_ _02849_ _02852_ _02850_ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__o21ai_1
XFILLER_50_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18329_ rbzero.spi_registers.got_new_other _02323_ _02283_ _02388_ vssd1 vssd1 vccd1
+ vccd1 _00833_ sky130_fd_sc_hd__a31o_1
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20222_ net282 _01153_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20153_ net213 _01084_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09964_ _03035_ vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20084_ clknet_leaf_84_i_clk _01015_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09895_ _02999_ vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10670_ _03462_ _03464_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__nor2_1
XFILLER_159_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12340_ _03487_ _05096_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__nand2_1
XFILLER_153_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12271_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[9\] vssd1
+ vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__or2_1
XFILLER_181_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19191__350 clknet_1_1__leaf__02750_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__inv_2
X_14010_ _06630_ _06752_ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__or2_1
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11222_ _02901_ _03838_ _03476_ _04006_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__a31o_1
X_19249__23 clknet_1_1__leaf__02755_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__inv_2
XFILLER_175_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11153_ rbzero.tex_r1\[56\] _03661_ _03936_ _03937_ vssd1 vssd1 vccd1 vccd1 _03938_
+ sky130_fd_sc_hd__a31o_1
XFILLER_122_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10104_ _03109_ vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__clkbuf_1
X_11084_ rbzero.map_overlay.i_otherx\[0\] _03462_ _03474_ rbzero.map_overlay.i_otherx\[3\]
+ _03869_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__a221o_1
X_15961_ _08524_ _08303_ vssd1 vssd1 vccd1 vccd1 _08577_ sky130_fd_sc_hd__and2_1
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10035_ _03072_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__clkbuf_4
X_14912_ _07585_ _07598_ vssd1 vssd1 vccd1 vccd1 _07600_ sky130_fd_sc_hd__and2_1
X_17700_ rbzero.debug_overlay.vplaneX\[0\] vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__buf_2
XFILLER_49_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18680_ _02411_ _02570_ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__nand2_1
X_15892_ _07693_ _07695_ _08509_ vssd1 vssd1 vccd1 vccd1 _08516_ sky130_fd_sc_hd__a21oi_1
XFILLER_91_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14843_ _06933_ _07048_ vssd1 vssd1 vccd1 vccd1 _07531_ sky130_fd_sc_hd__nor2_1
X_17631_ rbzero.debug_overlay.playerY\[4\] _03341_ _01908_ _01909_ vssd1 vssd1 vccd1
+ vccd1 _01910_ sky130_fd_sc_hd__a22o_1
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17562_ _01836_ _01839_ _01837_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__o21bai_1
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14774_ _07446_ _07460_ _07461_ vssd1 vssd1 vccd1 vccd1 _07462_ sky130_fd_sc_hd__a21oi_1
X_11986_ net47 _04730_ _04732_ _04759_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__a22o_1
XFILLER_189_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16513_ _09121_ _09122_ vssd1 vssd1 vccd1 vccd1 _09123_ sky130_fd_sc_hd__nor2_1
XFILLER_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19301_ rbzero.traced_texa\[-4\] rbzero.texV\[-4\] vssd1 vssd1 vccd1 vccd1 _02791_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_147_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13725_ _05527_ _05988_ _06480_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__o21bai_1
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10937_ rbzero.tex_r0\[45\] rbzero.tex_r0\[44\] _03690_ vssd1 vssd1 vccd1 vccd1 _03723_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17493_ _01784_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__clkbuf_4
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16444_ _09053_ _09054_ vssd1 vssd1 vccd1 vccd1 _09055_ sky130_fd_sc_hd__nor2_1
XFILLER_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13656_ _06370_ _06407_ _06412_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__and3_1
X_10868_ rbzero.tex_r0\[1\] rbzero.tex_r0\[0\] _03649_ vssd1 vssd1 vccd1 vccd1 _03654_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12607_ _05359_ _05363_ _05270_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__mux2_1
X_16375_ _08867_ _08869_ _08866_ vssd1 vssd1 vccd1 vccd1 _08986_ sky130_fd_sc_hd__a21bo_1
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13587_ _06001_ _06156_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__nor2_1
XFILLER_157_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ _03579_ _03584_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__nand2_1
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18114_ rbzero.spi_registers.new_other\[6\] _02264_ _02265_ _02266_ vssd1 vssd1 vccd1
+ vccd1 _00750_ sky130_fd_sc_hd__o211a_1
X_15326_ _07213_ _07757_ vssd1 vssd1 vccd1 vccd1 _08012_ sky130_fd_sc_hd__or2_1
XFILLER_184_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12538_ _05212_ _05256_ _05219_ _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__and4_1
XFILLER_158_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18045_ _02102_ _02103_ _02224_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__and3_1
X_15257_ _07856_ _07270_ _07855_ _07854_ vssd1 vssd1 vccd1 vccd1 _07943_ sky130_fd_sc_hd__o31ai_2
XFILLER_144_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12469_ _05198_ _05225_ _05207_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__or3b_2
XFILLER_67_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14208_ _06895_ _05096_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__mux2_1
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15188_ _07094_ _07732_ vssd1 vssd1 vccd1 vccd1 _07875_ sky130_fd_sc_hd__nand2_1
XFILLER_113_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14139_ _06834_ vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__clkbuf_1
X_19996_ clknet_leaf_94_i_clk _00927_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_140_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18878_ _04500_ _04499_ _02279_ _04507_ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a31o_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17829_ _02067_ _02077_ _02091_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__o21ai_1
XFILLER_39_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20205_ net265 _01136_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20136_ clknet_leaf_89_i_clk _01067_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
X_09947_ _03026_ vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20067_ clknet_3_4_0_i_clk _00998_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09878_ _02990_ vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__clkbuf_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ net12 net13 vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__nand2_1
XFILLER_79_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ net8 _04546_ _04547_ _04548_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__and4_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19254__4 clknet_1_0__leaf__02433_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__inv_2
XFILLER_14_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13510_ _06257_ _06266_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__xor2_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19223__379 clknet_1_0__leaf__02753_ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__inv_2
X_10722_ _03509_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__buf_4
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _07177_ vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__buf_2
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13441_ _06195_ _06197_ _06097_ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__a21o_1
X_10653_ _03446_ _03358_ rbzero.map_rom.a6 _03447_ _03448_ vssd1 vssd1 vccd1 vccd1
+ _03449_ sky130_fd_sc_hd__o221a_1
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16160_ _07494_ _08130_ vssd1 vssd1 vccd1 vccd1 _08773_ sky130_fd_sc_hd__or2_1
X_18390__34 clknet_1_1__leaf__02434_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__inv_2
XFILLER_127_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13372_ _06122_ _06128_ vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__nand2_1
XFILLER_107_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10584_ rbzero.debug_overlay.playerX\[0\] _03373_ rbzero.wall_tracer.mapX\[5\] _03378_
+ _03379_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__o221ai_1
XFILLER_10_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15111_ _07780_ _07798_ vssd1 vssd1 vccd1 vccd1 _07799_ sky130_fd_sc_hd__xnor2_4
X_12323_ _05062_ _05060_ _05072_ _05061_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__a211o_4
X_16091_ _08603_ _08704_ vssd1 vssd1 vccd1 vccd1 _08705_ sky130_fd_sc_hd__and2_1
XFILLER_182_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15042_ _07617_ _07137_ vssd1 vssd1 vccd1 vccd1 _07730_ sky130_fd_sc_hd__nor2_1
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12254_ _04926_ _04944_ _05013_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__and3_1
XFILLER_182_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11205_ rbzero.tex_r1\[18\] _03620_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__or2_1
XFILLER_134_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19850_ clknet_leaf_24_i_clk _00781_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_19117__284 clknet_1_1__leaf__02742_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__inv_2
X_12185_ rbzero.wall_tracer.state\[6\] vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__buf_4
X_18801_ rbzero.debug_overlay.facingY\[-3\] _02660_ vssd1 vssd1 vccd1 vccd1 _02661_
+ sky130_fd_sc_hd__or2_1
X_11136_ rbzero.tex_r1\[53\] _03652_ _03767_ _03673_ vssd1 vssd1 vccd1 vccd1 _03921_
+ sky130_fd_sc_hd__a31o_1
XFILLER_150_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19781_ clknet_leaf_81_i_clk _00712_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16993_ _09563_ _09598_ vssd1 vssd1 vccd1 vccd1 _09599_ sky130_fd_sc_hd__nand2_1
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18732_ rbzero.debug_overlay.playerY\[1\] _02582_ _02613_ _02559_ vssd1 vssd1 vccd1
+ vccd1 _01021_ sky130_fd_sc_hd__a211o_1
X_11067_ rbzero.map_overlay.i_mapdy\[2\] _03852_ gpout0.vpos\[7\] _03451_ vssd1 vssd1
+ vccd1 vccd1 _03853_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15944_ _08509_ vssd1 vssd1 vccd1 vccd1 _08562_ sky130_fd_sc_hd__clkbuf_4
XFILLER_114_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10018_ rbzero.tex_g1\[55\] rbzero.tex_g1\[56\] _03061_ vssd1 vssd1 vccd1 vccd1 _03064_
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18663_ rbzero.debug_overlay.playerX\[0\] _07032_ vssd1 vssd1 vccd1 vccd1 _02561_
+ sky130_fd_sc_hd__or2_1
XFILLER_49_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15875_ rbzero.wall_tracer.mapX\[9\] _07826_ _08498_ vssd1 vssd1 vccd1 vccd1 _08501_
+ sky130_fd_sc_hd__o21a_1
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18453__90 clknet_1_1__leaf__02441_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__inv_2
XFILLER_64_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17614_ _03390_ _04934_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__or2_1
X_14826_ _07456_ _07457_ vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__xnor2_1
X_18594_ _02516_ vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17545_ _01784_ rbzero.debug_overlay.vplaneY\[-3\] vssd1 vssd1 vccd1 vccd1 _01834_
+ sky130_fd_sc_hd__nor2_1
X_14757_ _07393_ _07406_ vssd1 vssd1 vccd1 vccd1 _07445_ sky130_fd_sc_hd__xnor2_1
X_11969_ net30 _04742_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__nor2_1
XFILLER_60_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13708_ _06450_ _06463_ _06464_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__a21o_1
X_17476_ _03340_ _01761_ _01767_ _01769_ vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__o22a_1
X_14688_ _07350_ _07352_ vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16427_ _09034_ _09037_ vssd1 vssd1 vccd1 vccd1 _09038_ sky130_fd_sc_hd__nand2_1
XFILLER_34_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13639_ _06349_ _06389_ _06390_ _06395_ vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__o31a_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16358_ _08858_ _08859_ _08856_ vssd1 vssd1 vccd1 vccd1 _08969_ sky130_fd_sc_hd__a21oi_1
XFILLER_118_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15309_ _07887_ _07890_ _07888_ vssd1 vssd1 vccd1 vccd1 _07995_ sky130_fd_sc_hd__o21ai_1
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16289_ _08898_ _08900_ vssd1 vssd1 vccd1 vccd1 _08901_ sky130_fd_sc_hd__nor2_1
XFILLER_161_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18028_ rbzero.pov.spi_buffer\[66\] rbzero.pov.ready_buffer\[66\] _02208_ vssd1 vssd1
+ vccd1 vccd1 _02216_ sky130_fd_sc_hd__mux2_1
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09801_ _02948_ vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19979_ net208 _00910_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09732_ _02912_ vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20119_ clknet_leaf_90_i_clk _01050_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_172_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13990_ _06588_ _06598_ _06605_ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__a21oi_1
XFILLER_58_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12941_ _05516_ _05471_ _05696_ _05697_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_58_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15660_ _08337_ _08338_ _08342_ vssd1 vssd1 vccd1 vccd1 _08343_ sky130_fd_sc_hd__a21oi_1
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12872_ _05604_ _05605_ _05627_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__or3_1
XFILLER_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _07297_ _07298_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__nand2_1
X_11823_ clknet_1_0__leaf__04486_ _04569_ _04577_ _04565_ _04599_ vssd1 vssd1 vccd1
+ vccd1 _04600_ sky130_fd_sc_hd__a32o_2
XFILLER_57_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _08273_ _08274_ vssd1 vssd1 vccd1 vccd1 _08275_ sky130_fd_sc_hd__xor2_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _01647_ _01648_ _01646_ vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__a21bo_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _07210_ _07228_ vssd1 vssd1 vccd1 vccd1 _07230_ sky130_fd_sc_hd__and2_1
XFILLER_187_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11754_ net52 vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__buf_4
XFILLER_121_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _01590_ _01591_ _01584_ _01587_ vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__a211oi_1
X_10705_ rbzero.wall_tracer.state\[1\] _03457_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__and2_1
XFILLER_41_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14473_ _06852_ _07160_ _03491_ vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__a21oi_4
X_11685_ _03689_ _04461_ _04465_ _03627_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__a211o_1
XFILLER_105_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16212_ _08823_ _08824_ vssd1 vssd1 vccd1 vccd1 _08825_ sky130_fd_sc_hd__and2b_1
XFILLER_128_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13424_ _06120_ _06133_ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__xnor2_1
X_10636_ _03430_ _03343_ _03352_ rbzero.map_overlay.i_othery\[0\] _03431_ vssd1 vssd1
+ vccd1 vccd1 _03432_ sky130_fd_sc_hd__a221o_1
X_17192_ rbzero.wall_tracer.trackDistY\[-10\] _01523_ _01533_ _08517_ vssd1 vssd1
+ vccd1 vccd1 _00561_ sky130_fd_sc_hd__o22a_1
XFILLER_139_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16143_ _08754_ _08755_ vssd1 vssd1 vccd1 vccd1 _08756_ sky130_fd_sc_hd__nor2_1
XFILLER_6_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13355_ _06103_ _06056_ _06111_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__o21a_1
XFILLER_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10567_ rbzero.debug_overlay.playerX\[2\] vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__inv_2
XFILLER_154_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12306_ _05061_ _05062_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__or2b_1
X_16074_ _08403_ _08405_ vssd1 vssd1 vccd1 vccd1 _08688_ sky130_fd_sc_hd__nand2_1
X_13286_ _05965_ _06018_ _06017_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__o21ba_1
X_10498_ rbzero.tex_b0\[20\] rbzero.tex_b0\[19\] _03313_ vssd1 vssd1 vccd1 vccd1 _03316_
+ sky130_fd_sc_hd__mux2_1
XFILLER_142_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15025_ _06900_ _07037_ vssd1 vssd1 vccd1 vccd1 _07713_ sky130_fd_sc_hd__or2_1
X_19902_ clknet_leaf_19_i_clk _00833_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_other
+ sky130_fd_sc_hd__dfxtp_1
X_12237_ _04958_ rbzero.wall_tracer.trackDistX\[6\] rbzero.wall_tracer.trackDistX\[5\]
+ _04959_ _04998_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__a221o_1
XFILLER_123_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19833_ clknet_leaf_4_i_clk _00764_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12168_ _03359_ _03351_ _04929_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__a21oi_1
XFILLER_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11119_ _03519_ _03900_ _03901_ _03903_ _03904_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__a41o_1
X_19764_ clknet_leaf_85_i_clk _00695_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_16976_ _09142_ _09231_ _09229_ _09133_ vssd1 vssd1 vccd1 vccd1 _09582_ sky130_fd_sc_hd__o22ai_1
X_12099_ rbzero.debug_overlay.facingY\[-8\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__nand2_1
XFILLER_83_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18715_ _06982_ _02535_ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__nor2_1
Xinput6 i_gpout0_sel[3] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_6
X_15927_ rbzero.wall_tracer.trackDistX\[-6\] rbzero.wall_tracer.stepDistX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _08547_ sky130_fd_sc_hd__or2_1
X_19695_ clknet_leaf_75_i_clk _00626_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18646_ rbzero.pov.ready_buffer\[63\] _06946_ _02540_ vssd1 vssd1 vccd1 vccd1 _02549_
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15858_ _08485_ _08487_ vssd1 vssd1 vccd1 vccd1 _08488_ sky130_fd_sc_hd__nor2_2
XFILLER_40_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14809_ _07487_ _07493_ _07496_ vssd1 vssd1 vccd1 vccd1 _07497_ sky130_fd_sc_hd__a21oi_2
X_18577_ _02507_ vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__clkbuf_1
X_15789_ _08448_ vssd1 vssd1 vccd1 vccd1 _08456_ sky130_fd_sc_hd__clkbuf_4
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17528_ _01757_ rbzero.debug_overlay.vplaneY\[-4\] vssd1 vssd1 vccd1 vccd1 _01818_
+ sky130_fd_sc_hd__or2_1
XFILLER_71_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17459_ rbzero.debug_overlay.vplaneY\[-5\] _01753_ vssd1 vssd1 vccd1 vccd1 _01754_
+ sky130_fd_sc_hd__xor2_1
XFILLER_178_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20470_ net126 _01401_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11470_ rbzero.tex_g1\[25\] rbzero.tex_g1\[24\] _04247_ vssd1 vssd1 vccd1 vccd1 _04253_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10421_ _03275_ vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ _05687_ _05761_ _05763_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__or3_1
X_10352_ _03239_ vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19034__208 clknet_1_1__leaf__02735_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__inv_2
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13071_ _05802_ _05824_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__xnor2_1
X_10283_ _03203_ vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12022_ net43 _04794_ net35 net36 vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__a211o_1
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16830_ _09435_ _09436_ vssd1 vssd1 vccd1 vccd1 _09437_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16761_ _09366_ _09367_ vssd1 vssd1 vccd1 vccd1 _09369_ sky130_fd_sc_hd__and2_1
XFILLER_150_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13973_ _05270_ _06652_ _06629_ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__a21o_1
XFILLER_24_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18500_ _02467_ vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15712_ _08389_ _08394_ vssd1 vssd1 vccd1 vccd1 _08395_ sky130_fd_sc_hd__xnor2_2
X_12924_ _05653_ _05660_ _05663_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__nor3_1
X_16692_ _09095_ _09300_ vssd1 vssd1 vccd1 vccd1 _09301_ sky130_fd_sc_hd__xnor2_1
X_19229__385 clknet_1_0__leaf__02753_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__inv_2
X_19480_ clknet_leaf_49_i_clk _00426_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_19_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15643_ _07972_ _08081_ _07959_ _07856_ vssd1 vssd1 vccd1 vccd1 _08326_ sky130_fd_sc_hd__o22a_1
XFILLER_132_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12855_ _05608_ _05611_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__xnor2_1
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _04565_ _04574_ _04582_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__a21o_1
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15574_ _08256_ _08257_ vssd1 vssd1 vccd1 vccd1 _08258_ sky130_fd_sc_hd__and2_1
X_18362_ rbzero.pov.spi_counter\[2\] rbzero.pov.spi_counter\[1\] rbzero.pov.spi_counter\[0\]
+ _02419_ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__and4bb_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12786_ _05541_ _05542_ _05355_ _05425_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17313_ _01636_ _01637_ vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__xnor2_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _07148_ vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__clkbuf_4
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ net4 net3 vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__and2_1
XFILLER_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18293_ rbzero.spi_registers.spi_buffer\[0\] rbzero.spi_registers.new_leak\[0\] _02379_
+ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__mux2_1
XFILLER_186_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14456_ _04947_ _06859_ vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__nor2_1
X_17244_ rbzero.wall_tracer.trackDistY\[-2\] rbzero.wall_tracer.stepDistY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__or2_1
X_11668_ _03607_ _04444_ _04448_ _03627_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__a211o_1
XFILLER_186_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13407_ _06162_ _06163_ vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__or2b_1
XFILLER_179_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17175_ _01516_ _01517_ _01515_ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__a21oi_1
X_10619_ _03413_ _03374_ rbzero.map_rom.a6 _03353_ _03414_ vssd1 vssd1 vccd1 vccd1
+ _03415_ sky130_fd_sc_hd__a221o_1
XFILLER_128_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14387_ _07010_ _07063_ _07074_ vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__a21oi_1
X_11599_ _04379_ _04380_ _03739_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__mux2_1
XFILLER_31_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16126_ _08737_ _08738_ vssd1 vssd1 vccd1 vccd1 _08739_ sky130_fd_sc_hd__nand2_1
XFILLER_6_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13338_ _06085_ _06094_ vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__xor2_1
XFILLER_182_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16057_ _08661_ _08670_ vssd1 vssd1 vccd1 vccd1 _08671_ sky130_fd_sc_hd__xnor2_2
XFILLER_143_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13269_ _05927_ _05969_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__nor2_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15008_ _07572_ _07610_ _07693_ _07695_ vssd1 vssd1 vccd1 vccd1 _07696_ sky130_fd_sc_hd__a22o_2
XFILLER_97_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19816_ clknet_leaf_1_i_clk _00747_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19747_ clknet_leaf_92_i_clk _00678_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16959_ _09498_ _09477_ vssd1 vssd1 vccd1 vccd1 _09565_ sky130_fd_sc_hd__or2b_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19678_ clknet_leaf_80_i_clk _00609_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18629_ _07145_ rbzero.pov.ready_buffer\[59\] _02535_ vssd1 vssd1 vccd1 vccd1 _02536_
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_3_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_11 _06855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_22 rbzero.spi_registers.vshift\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_33 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20522_ clknet_leaf_41_i_clk _01453_ vssd1 vssd1 vccd1 vccd1 gpout3.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_44 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_55 _01786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_66 net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20453_ net133 _01384_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20384_ net444 _01315_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10970_ rbzero.tex_r0\[55\] rbzero.tex_r0\[54\] _03690_ vssd1 vssd1 vccd1 vccd1 _03756_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12640_ _05269_ _05329_ _05378_ _05384_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__and4_1
XFILLER_93_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12571_ _05310_ _05316_ _05323_ _05327_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__o211a_1
XFILLER_62_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14310_ _06966_ _06977_ vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__or2_1
X_11522_ _04198_ _04300_ _04304_ _03721_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__a211o_1
XFILLER_54_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15290_ _07972_ _07270_ _07975_ vssd1 vssd1 vccd1 vccd1 _07976_ sky130_fd_sc_hd__or3_1
XFILLER_141_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14241_ _06927_ _06928_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__nand2_1
XFILLER_172_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11453_ _03540_ _03632_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__nor2_2
XFILLER_183_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10404_ _03266_ vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14172_ _06859_ vssd1 vssd1 vccd1 vccd1 _06860_ sky130_fd_sc_hd__buf_2
X_11384_ _03674_ _04163_ _04167_ _03679_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__a211o_1
XFILLER_152_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13123_ _05879_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__dlymetal6s2s_1
X_10335_ _03230_ vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13054_ _05488_ _05810_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__xnor2_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17931_ _02165_ vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__clkbuf_1
X_10266_ _03194_ vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12005_ _04393_ _04723_ _04726_ _04770_ _04778_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__a32oi_2
XFILLER_120_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17862_ rbzero.spi_registers.sclk_buffer\[2\] rbzero.spi_registers.sclk_buffer\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__nand2b_2
X_10197_ _03158_ vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19601_ clknet_leaf_31_i_clk _00532_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.wall\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_16813_ _09417_ _09418_ _09419_ vssd1 vssd1 vccd1 vccd1 _09421_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17793_ _02046_ _02047_ _02045_ vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__a21o_1
XFILLER_94_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19532_ clknet_leaf_58_i_clk _00004_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_16744_ _09264_ _09323_ _09350_ vssd1 vssd1 vccd1 vccd1 _09352_ sky130_fd_sc_hd__nand3_1
X_13956_ rbzero.wall_tracer.stepDistY\[-4\] _06705_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _06706_ sky130_fd_sc_hd__mux2_1
XFILLER_35_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12907_ _05653_ _05660_ _05663_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__o21a_1
XFILLER_35_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19463_ clknet_leaf_56_i_clk _00409_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16675_ _09279_ _09283_ vssd1 vssd1 vccd1 vccd1 _09284_ sky130_fd_sc_hd__xnor2_1
XFILLER_59_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13887_ _06640_ _06642_ _06603_ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__mux2_1
XFILLER_185_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18945__128 clknet_1_0__leaf__02726_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__inv_2
X_12838_ _05591_ _05594_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__nor2_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15626_ _08182_ _08308_ _04832_ vssd1 vssd1 vccd1 vccd1 _08310_ sky130_fd_sc_hd__a21o_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19394_ rbzero.traced_texVinit\[1\] _08463_ _07813_ _08455_ vssd1 vssd1 vccd1 vccd1
+ _01429_ sky130_fd_sc_hd__a22o_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18345_ rbzero.spi_registers.got_new_vshift _02323_ _02283_ _02401_ vssd1 vssd1 vccd1
+ vccd1 _00840_ sky130_fd_sc_hd__a31o_1
X_15557_ _08125_ _08223_ _08239_ vssd1 vssd1 vccd1 vccd1 _08241_ sky130_fd_sc_hd__nand3_1
X_12769_ _05210_ _05424_ _05417_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__nand3_4
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14508_ _07195_ _04948_ _03492_ _07134_ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__nor4_2
XFILLER_174_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15488_ _08064_ _08172_ vssd1 vssd1 vccd1 vccd1 _08173_ sky130_fd_sc_hd__xnor2_2
X_18276_ _02369_ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__clkbuf_4
XFILLER_175_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput20 i_gpout2_sel[5] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_4
X_17227_ _01560_ _01561_ _01562_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__o21ai_1
XFILLER_174_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput31 i_gpout4_sel[4] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_4
X_14439_ _07125_ _07126_ vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__nand2_1
XFILLER_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput42 i_reg_csb vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_8
Xinput53 i_vec_sclk vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_8
XFILLER_116_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17158_ _01499_ _01501_ vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__xnor2_1
XFILLER_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16109_ _08635_ _08604_ vssd1 vssd1 vccd1 vccd1 _08722_ sky130_fd_sc_hd__or2b_1
X_09980_ rbzero.tex_r0\[10\] rbzero.tex_r0\[9\] _03039_ vssd1 vssd1 vccd1 vccd1 _03044_
+ sky130_fd_sc_hd__mux2_1
X_17089_ _09597_ _09564_ vssd1 vssd1 vccd1 vccd1 _09694_ sky130_fd_sc_hd__and2b_1
Xclkbuf_1_1__f__02747_ clknet_0__02747_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02747_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_170_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20505_ clknet_leaf_42_i_clk _01436_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19232__7 clknet_1_1__leaf__02754_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__inv_2
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20436_ net496 _01367_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20367_ net427 _01298_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[22\] sky130_fd_sc_hd__dfxtp_1
X_10120_ rbzero.tex_g1\[7\] rbzero.tex_g1\[8\] _03117_ vssd1 vssd1 vccd1 vccd1 _03118_
+ sky130_fd_sc_hd__mux2_1
XFILLER_121_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20298_ net358 _01229_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[17\] sky130_fd_sc_hd__dfxtp_1
X_10051_ _03081_ vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19146__309 clknet_1_1__leaf__02746_ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__inv_2
XFILLER_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13810_ _06280_ _06330_ _06331_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__and3_1
X_14790_ _07471_ _07477_ vssd1 vssd1 vccd1 vccd1 _07478_ sky130_fd_sc_hd__nand2_1
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13741_ _05503_ _06230_ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__or2_1
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10953_ _03635_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__buf_6
XFILLER_189_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16460_ _08972_ _09070_ vssd1 vssd1 vccd1 vccd1 _09071_ sky130_fd_sc_hd__xnor2_2
X_13672_ _06354_ _06381_ _06428_ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__a21oi_1
X_10884_ _03669_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__buf_4
XFILLER_25_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15411_ _08095_ _08004_ vssd1 vssd1 vccd1 vccd1 _08096_ sky130_fd_sc_hd__nand2_1
X_12623_ _05330_ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__clkbuf_4
X_16391_ _08905_ _08974_ _09001_ vssd1 vssd1 vccd1 vccd1 _09002_ sky130_fd_sc_hd__a21o_1
XFILLER_58_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15342_ _08026_ _08027_ vssd1 vssd1 vccd1 vccd1 _08028_ sky130_fd_sc_hd__nand2_1
X_18130_ rbzero.spi_registers.new_other\[2\] _02264_ _02274_ _02275_ vssd1 vssd1 vccd1
+ vccd1 _00757_ sky130_fd_sc_hd__o211a_1
XFILLER_169_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12554_ _05307_ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__clkbuf_4
XFILLER_185_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11505_ _04198_ _04287_ _03721_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__a21o_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15273_ rbzero.wall_tracer.visualWallDist\[7\] _07256_ vssd1 vssd1 vccd1 vccd1 _07959_
+ sky130_fd_sc_hd__nand2_2
XFILLER_129_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18061_ _02234_ vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__clkbuf_1
X_12485_ _05114_ _05241_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__xnor2_4
XFILLER_185_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17012_ _09617_ _09516_ _09515_ vssd1 vssd1 vccd1 vccd1 _09618_ sky130_fd_sc_hd__a21o_1
XFILLER_156_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14224_ rbzero.debug_overlay.playerX\[-8\] rbzero.debug_overlay.playerX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__xnor2_1
X_11436_ rbzero.tex_g0\[42\] _03649_ _03610_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__a21o_1
XFILLER_144_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14155_ _06845_ vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__clkbuf_1
X_11367_ rbzero.tex_g0\[21\] rbzero.tex_g0\[20\] _03709_ vssd1 vssd1 vccd1 vccd1 _04151_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13106_ _05301_ _05862_ _05610_ _05355_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__o22a_1
X_10318_ rbzero.tex_b1\[41\] rbzero.tex_b1\[42\] _03221_ vssd1 vssd1 vccd1 vccd1 _03222_
+ sky130_fd_sc_hd__mux2_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14086_ rbzero.wall_tracer.trackDistX\[3\] _06788_ _06806_ vssd1 vssd1 vccd1 vccd1
+ _00442_ sky130_fd_sc_hd__o21a_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _04065_ _04082_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__nor2_4
XFILLER_79_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _05791_ _05793_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__or2_1
X_17914_ _02156_ vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__clkbuf_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10249_ _03185_ vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18894_ _03515_ _02714_ _02323_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__o21a_1
XFILLER_6_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17845_ rbzero.spi_registers.spi_counter\[3\] rbzero.spi_registers.spi_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__or2_1
XFILLER_66_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19012__188 clknet_1_1__leaf__02733_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__inv_2
XFILLER_94_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19086__256 clknet_1_1__leaf__02739_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__inv_2
X_17776_ _01985_ rbzero.debug_overlay.vplaneX\[-3\] vssd1 vssd1 vccd1 vccd1 _02043_
+ sky130_fd_sc_hd__and2_1
XFILLER_94_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14988_ _07671_ _07674_ _07668_ vssd1 vssd1 vccd1 vccd1 _07676_ sky130_fd_sc_hd__o21ai_1
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19515_ clknet_leaf_52_i_clk _00461_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16727_ _08888_ _09110_ _09234_ _09233_ vssd1 vssd1 vccd1 vccd1 _09335_ sky130_fd_sc_hd__o31ai_2
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13939_ _06618_ _06624_ vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__nor2_1
XFILLER_74_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19446_ _02334_ _02893_ _02894_ vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__and3_1
X_16658_ _09246_ _09266_ vssd1 vssd1 vccd1 vccd1 _09267_ sky130_fd_sc_hd__xnor2_2
XFILLER_62_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_83_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_15609_ _08187_ _08292_ vssd1 vssd1 vccd1 vccd1 _08293_ sky130_fd_sc_hd__xnor2_1
X_19377_ rbzero.traced_texa\[8\] rbzero.texV\[8\] vssd1 vssd1 vccd1 vccd1 _02855_
+ sky130_fd_sc_hd__nand2_1
X_16589_ rbzero.wall_tracer.trackDistX\[4\] rbzero.wall_tracer.stepDistX\[4\] vssd1
+ vssd1 vccd1 vccd1 _09199_ sky130_fd_sc_hd__or2_1
XFILLER_188_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18328_ _02398_ vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__clkbuf_1
XFILLER_187_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18259_ _02107_ rbzero.spi_registers.spi_cmd\[1\] _02981_ _02359_ vssd1 vssd1 vccd1
+ vccd1 _02360_ sky130_fd_sc_hd__or4_1
XFILLER_128_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20221_ net281 _01152_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_21_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_09963_ rbzero.tex_r0\[18\] rbzero.tex_r0\[17\] _03028_ vssd1 vssd1 vccd1 vccd1 _03035_
+ sky130_fd_sc_hd__mux2_1
X_20152_ clknet_leaf_18_i_clk _01083_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_mapd
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09894_ rbzero.tex_r0\[51\] rbzero.tex_r0\[50\] _02995_ vssd1 vssd1 vccd1 vccd1 _02999_
+ sky130_fd_sc_hd__mux2_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20083_ clknet_leaf_84_i_clk _01014_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_100_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12270_ _05007_ _05026_ _05027_ _05009_ rbzero.wall_tracer.mapY\[10\] vssd1 vssd1
+ vccd1 vccd1 _00405_ sky130_fd_sc_hd__a32o_1
XFILLER_135_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11221_ _03460_ _03467_ _03525_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__nor3_1
XFILLER_88_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20419_ net479 _01350_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11152_ rbzero.tex_r1\[57\] _03919_ _03768_ _03670_ vssd1 vssd1 vccd1 vccd1 _03937_
+ sky130_fd_sc_hd__a31o_1
XFILLER_136_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10103_ rbzero.tex_g1\[15\] rbzero.tex_g1\[16\] _03106_ vssd1 vssd1 vccd1 vccd1 _03109_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11083_ rbzero.map_overlay.i_otherx\[4\] _02900_ vssd1 vssd1 vccd1 vccd1 _03869_
+ sky130_fd_sc_hd__xor2_1
X_15960_ _08569_ _08489_ _08576_ vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__a21oi_1
XFILLER_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10034_ _02908_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__buf_4
X_14911_ _07585_ _07598_ vssd1 vssd1 vccd1 vccd1 _07599_ sky130_fd_sc_hd__nor2_1
XFILLER_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15891_ rbzero.wall_tracer.trackDistX\[-11\] _08508_ _08511_ _08515_ vssd1 vssd1
+ vccd1 vccd1 _00538_ sky130_fd_sc_hd__o22a_1
XFILLER_48_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17630_ _03341_ _04943_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__nor2_1
X_14842_ _06970_ vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__clkbuf_4
XFILLER_36_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17561_ _01847_ _01848_ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__nand2_1
XFILLER_91_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11985_ net52 _04723_ net48 vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__a21o_1
X_14773_ _07447_ _07459_ vssd1 vssd1 vccd1 vccd1 _07461_ sky130_fd_sc_hd__and2b_1
XFILLER_189_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19300_ _02759_ _02789_ _02790_ _02762_ rbzero.texV\[-5\] vssd1 vssd1 vccd1 vccd1
+ _01412_ sky130_fd_sc_hd__a32o_1
X_16512_ _08986_ _08995_ _08993_ vssd1 vssd1 vccd1 vccd1 _09122_ sky130_fd_sc_hd__a21oi_1
XFILLER_56_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10936_ rbzero.tex_r0\[47\] rbzero.tex_r0\[46\] _03664_ vssd1 vssd1 vccd1 vccd1 _03722_
+ sky130_fd_sc_hd__mux2_1
X_13724_ _05527_ _05987_ _06480_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__or3b_1
XFILLER_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17492_ rbzero.debug_overlay.vplaneY\[10\] vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__buf_2
XFILLER_140_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19231_ clknet_1_1__leaf__04486_ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__buf_1
XFILLER_108_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16443_ _08807_ _08926_ _08805_ vssd1 vssd1 vccd1 vccd1 _09054_ sky130_fd_sc_hd__a21boi_1
XFILLER_147_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10867_ _03650_ _03651_ _03652_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__mux2_1
X_13655_ _06368_ _06408_ _06409_ _06411_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__a22o_1
XFILLER_182_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12606_ _05361_ _05362_ _05338_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__mux2_1
X_16374_ _08983_ _08984_ vssd1 vssd1 vccd1 vccd1 _08985_ sky130_fd_sc_hd__xor2_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ _06341_ _06336_ vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__xor2_1
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _03577_ _03578_ rbzero.texV\[7\] vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__a21o_1
XFILLER_185_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19200__358 clknet_1_0__leaf__02751_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__inv_2
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18113_ _04828_ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__clkbuf_4
X_15325_ _08007_ _08010_ vssd1 vssd1 vccd1 vccd1 _08011_ sky130_fd_sc_hd__xnor2_1
X_12537_ _05217_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__inv_2
XFILLER_185_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18044_ rbzero.spi_registers.spi_counter\[6\] rbzero.spi_registers.spi_counter\[5\]
+ rbzero.spi_registers.spi_counter\[4\] _02106_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__or4_1
XFILLER_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15256_ _07873_ _07851_ vssd1 vssd1 vccd1 vccd1 _07942_ sky130_fd_sc_hd__or2b_1
X_12468_ _05146_ _05200_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__xnor2_2
XFILLER_138_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11419_ rbzero.tex_g0\[63\] rbzero.tex_g0\[62\] _03699_ vssd1 vssd1 vccd1 vccd1 _04203_
+ sky130_fd_sc_hd__mux2_1
XFILLER_160_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14207_ _04904_ vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__clkinv_2
X_15187_ _07851_ _07873_ vssd1 vssd1 vccd1 vccd1 _07874_ sky130_fd_sc_hd__xnor2_1
X_12399_ rbzero.wall_tracer.visualWallDist\[5\] _03480_ vssd1 vssd1 vccd1 vccd1 _05156_
+ sky130_fd_sc_hd__nor2_1
XFILLER_153_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14138_ rbzero.wall_tracer.stepDistX\[6\] _06767_ _06825_ vssd1 vssd1 vccd1 vccd1
+ _06834_ sky130_fd_sc_hd__mux2_1
XFILLER_193_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19995_ clknet_leaf_94_i_clk _00926_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14069_ rbzero.wall_tracer.visualWallDist\[-5\] _06796_ _06785_ rbzero.wall_tracer.trackDistY\[-5\]
+ _06797_ vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__o221a_1
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18877_ _04500_ _02286_ _02705_ _02285_ vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__o211a_1
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17828_ rbzero.wall_tracer.rayAddendX\[8\] rbzero.wall_tracer.rayAddendX\[7\] _02001_
+ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__o21ai_1
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17759_ _02018_ _02023_ _02026_ vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__o21a_1
XFILLER_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19429_ rbzero.wall_tracer.rayAddendX\[-7\] _08448_ _08454_ _02884_ vssd1 vssd1 vccd1
+ vccd1 _01447_ sky130_fd_sc_hd__a22o_1
XFILLER_62_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18997__176 clknet_1_1__leaf__02730_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__inv_2
XFILLER_159_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20204_ net264 _01135_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20135_ clknet_leaf_78_i_clk _01066_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
X_09946_ rbzero.tex_r0\[26\] rbzero.tex_r0\[25\] _03017_ vssd1 vssd1 vccd1 vccd1 _03026_
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20066_ clknet_leaf_83_i_clk _00997_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_100_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09877_ rbzero.tex_r0\[59\] rbzero.tex_r0\[58\] _02984_ vssd1 vssd1 vccd1 vccd1 _02990_
+ sky130_fd_sc_hd__mux2_1
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19069__240 clknet_1_0__leaf__02738_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__inv_2
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ net6 _04496_ net7 vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__a21o_1
XFILLER_198_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10721_ _03508_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__clkinv_4
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _06104_ _06107_ _06196_ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__a21o_1
XFILLER_201_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10652_ rbzero.map_overlay.i_mapdy\[2\] rbzero.map_rom.b6 vssd1 vssd1 vccd1 vccd1
+ _03448_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13371_ _06002_ _06034_ _06054_ _06121_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__a211o_1
X_10583_ _03378_ rbzero.wall_tracer.mapX\[5\] rbzero.wall_tracer.mapX\[7\] rbzero.wall_tracer.mapX\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__a211oi_1
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15110_ _07796_ _07797_ vssd1 vssd1 vccd1 vccd1 _07798_ sky130_fd_sc_hd__nor2_2
X_12322_ rbzero.wall_tracer.visualWallDist\[4\] _03480_ vssd1 vssd1 vccd1 vccd1 _05079_
+ sky130_fd_sc_hd__nor2_1
X_16090_ _08702_ _08703_ vssd1 vssd1 vccd1 vccd1 _08704_ sky130_fd_sc_hd__xor2_1
XFILLER_6_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15041_ _07110_ vssd1 vssd1 vccd1 vccd1 _07729_ sky130_fd_sc_hd__inv_2
XFILLER_170_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12253_ _05010_ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__clkinv_2
XFILLER_108_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11204_ rbzero.tex_r1\[20\] _03920_ _03936_ _03987_ _03988_ vssd1 vssd1 vccd1 vccd1
+ _03989_ sky130_fd_sc_hd__a311o_1
XFILLER_141_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12184_ _03341_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__buf_4
XFILLER_69_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18800_ _02637_ vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__clkbuf_2
X_11135_ _03919_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__clkbuf_4
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19780_ clknet_leaf_81_i_clk _00711_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_16992_ _09564_ _09597_ vssd1 vssd1 vccd1 vccd1 _09598_ sky130_fd_sc_hd__xnor2_1
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18731_ rbzero.pov.ready_buffer\[54\] _02411_ _02535_ _02612_ _02587_ vssd1 vssd1
+ vccd1 vccd1 _02613_ sky130_fd_sc_hd__o221a_1
XFILLER_77_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11066_ _03849_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__buf_4
X_15943_ _08524_ _08052_ vssd1 vssd1 vccd1 vccd1 _08561_ sky130_fd_sc_hd__and2_1
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10017_ _03063_ vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__clkbuf_1
X_18662_ rbzero.debug_overlay.playerX\[0\] _07032_ vssd1 vssd1 vccd1 vccd1 _02560_
+ sky130_fd_sc_hd__nand2_1
XFILLER_95_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ rbzero.wall_tracer.mapX\[9\] _08489_ _08488_ _08500_ vssd1 vssd1 vccd1 vccd1
+ _00536_ sky130_fd_sc_hd__a22o_1
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17613_ _01895_ vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14825_ _07492_ _07488_ vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__xnor2_1
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18593_ rbzero.pov.spi_buffer\[64\] rbzero.pov.spi_buffer\[65\] _02510_ vssd1 vssd1
+ vccd1 vccd1 _02516_ sky130_fd_sc_hd__mux2_1
XFILLER_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17544_ _01830_ _01831_ _01829_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__a21o_1
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14756_ _07409_ _07422_ vssd1 vssd1 vccd1 vccd1 _07444_ sky130_fd_sc_hd__xnor2_1
X_11968_ net29 vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__inv_2
XFILLER_45_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13707_ _06451_ _06462_ vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__and2_1
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10919_ _03689_ _03694_ _03703_ _03704_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__a211o_1
XFILLER_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17475_ _03339_ _01768_ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__nand2_1
X_11899_ _02899_ _03527_ _03526_ _04020_ net21 net22 vssd1 vssd1 vccd1 vccd1 _04674_
+ sky130_fd_sc_hd__mux4_1
X_14687_ _07355_ _07356_ vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__xnor2_1
X_19124__289 clknet_1_0__leaf__02744_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__inv_2
XFILLER_189_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16426_ _08245_ _09035_ _09036_ _08247_ vssd1 vssd1 vccd1 vccd1 _09037_ sky130_fd_sc_hd__o22ai_1
X_13638_ _06392_ _06394_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__nand2_1
XFILLER_34_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16357_ _08881_ _08847_ vssd1 vssd1 vccd1 vccd1 _08968_ sky130_fd_sc_hd__or2b_1
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13569_ _06307_ _06324_ _06325_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__a21oi_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15308_ _07992_ _07993_ _07882_ vssd1 vssd1 vccd1 vccd1 _07994_ sky130_fd_sc_hd__or3_1
XFILLER_173_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19076_ clknet_1_0__leaf__02732_ vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__buf_1
X_16288_ _08108_ _08899_ _08775_ _08774_ vssd1 vssd1 vccd1 vccd1 _08900_ sky130_fd_sc_hd__o31a_1
XFILLER_117_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18027_ _02215_ vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15239_ _07336_ _07802_ _07925_ vssd1 vssd1 vccd1 vccd1 _07926_ sky130_fd_sc_hd__a21oi_2
XFILLER_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09800_ rbzero.tex_r1\[29\] rbzero.tex_r1\[30\] _02943_ vssd1 vssd1 vccd1 vccd1 _02948_
+ sky130_fd_sc_hd__mux2_1
X_19018__194 clknet_1_0__leaf__02733_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__inv_2
XFILLER_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19978_ net207 _00909_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09731_ rbzero.tex_r1\[62\] rbzero.tex_r1\[63\] _02910_ vssd1 vssd1 vccd1 vccd1 _02912_
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20118_ clknet_leaf_90_i_clk _01049_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
X_09929_ _02983_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__clkbuf_4
XFILLER_172_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20049_ clknet_leaf_82_i_clk _00980_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[65\]
+ sky130_fd_sc_hd__dfxtp_1
X_12940_ _05534_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__clkbuf_4
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _05604_ _05605_ _05627_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__o21ai_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _07092_ _07147_ vssd1 vssd1 vccd1 vccd1 _07298_ sky130_fd_sc_hd__nor2_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ net53 _04569_ _04568_ net51 _04598_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__a221o_1
X_15590_ _08138_ _08146_ _08143_ vssd1 vssd1 vccd1 vccd1 _08274_ sky130_fd_sc_hd__a21bo_1
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _04496_ _04530_ net6 vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__and3b_1
X_14541_ _07210_ _07228_ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__nor2_1
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _03492_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__buf_4
XFILLER_186_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17260_ _01584_ _01587_ _01590_ _01591_ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__o211a_1
XFILLER_198_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11684_ _03656_ _04462_ _04463_ _04464_ _03673_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__o221a_1
X_14472_ _04881_ _05171_ _06849_ vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__mux2_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16211_ _08821_ _08822_ vssd1 vssd1 vccd1 vccd1 _08824_ sky130_fd_sc_hd__nand2_1
X_13423_ _06177_ _06179_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__nand2_1
X_10635_ rbzero.map_overlay.i_otherx\[3\] _03369_ vssd1 vssd1 vccd1 vccd1 _03431_
+ sky130_fd_sc_hd__xor2_1
X_17191_ _08562_ _01531_ _01532_ _01527_ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__a31o_1
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16142_ _08617_ _08626_ _08624_ vssd1 vssd1 vccd1 vccd1 _08755_ sky130_fd_sc_hd__a21oi_1
XFILLER_10_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13354_ _06104_ _06105_ _06109_ _06110_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__a31o_1
X_10566_ _03343_ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__clkinv_2
XFILLER_127_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12305_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[10\] vssd1
+ vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__nand2_1
XFILLER_155_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16073_ _08676_ _08686_ vssd1 vssd1 vccd1 vccd1 _08687_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13285_ _06011_ _06041_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__xnor2_1
X_10497_ _03315_ vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15024_ _07710_ _07711_ vssd1 vssd1 vccd1 vccd1 _07712_ sky130_fd_sc_hd__xnor2_1
X_19901_ clknet_leaf_15_i_clk _00832_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_12236_ rbzero.wall_tracer.trackDistX\[5\] _04959_ _04960_ rbzero.wall_tracer.trackDistX\[4\]
+ _04997_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__o221a_1
XFILLER_170_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19832_ clknet_leaf_4_i_clk _00763_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12167_ _04928_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__clkbuf_4
XFILLER_111_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11118_ _03502_ _03518_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__nand2_1
XFILLER_1_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19763_ clknet_leaf_85_i_clk _00694_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_16975_ _09133_ _09142_ _09231_ _09229_ vssd1 vssd1 vccd1 vccd1 _09581_ sky130_fd_sc_hd__or4_1
X_12098_ rbzero.debug_overlay.facingY\[-8\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18714_ rbzero.debug_overlay.playerY\[-4\] _02588_ _02600_ _02586_ vssd1 vssd1 vccd1
+ vccd1 _01016_ sky130_fd_sc_hd__o211a_1
XFILLER_77_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11049_ _03834_ rbzero.debug_overlay.playerY\[1\] vssd1 vssd1 vccd1 vccd1 _03835_
+ sky130_fd_sc_hd__xnor2_1
X_15926_ _08524_ _07808_ vssd1 vssd1 vccd1 vccd1 _08546_ sky130_fd_sc_hd__and2_1
X_19694_ clknet_leaf_9_i_clk _00625_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[5\]
+ sky130_fd_sc_hd__dfxtp_2
Xinput7 i_gpout0_sel[4] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_6
X_18645_ _02534_ _02547_ _02548_ _02356_ vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__o211a_1
XFILLER_92_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ _08486_ vssd1 vssd1 vccd1 vccd1 _08487_ sky130_fd_sc_hd__buf_2
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14808_ _07411_ _07495_ vssd1 vssd1 vccd1 vccd1 _07496_ sky130_fd_sc_hd__or2_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18576_ rbzero.pov.spi_buffer\[56\] rbzero.pov.spi_buffer\[57\] _02499_ vssd1 vssd1
+ vccd1 vccd1 _02507_ sky130_fd_sc_hd__mux2_1
XFILLER_80_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15788_ rbzero.row_render.size\[3\] _08449_ _06695_ _08455_ vssd1 vssd1 vccd1 vccd1
+ _00495_ sky130_fd_sc_hd__a22o_1
XFILLER_45_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19206__364 clknet_1_1__leaf__02751_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__inv_2
X_17527_ _01814_ _01801_ _01815_ _03339_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__a31o_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14739_ _07425_ _07426_ vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__xnor2_2
XFILLER_178_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17458_ rbzero.debug_overlay.vplaneY\[-6\] rbzero.debug_overlay.vplaneY\[-7\] rbzero.debug_overlay.vplaneY\[-8\]
+ _01752_ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__o31a_1
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16409_ _09018_ _09019_ vssd1 vssd1 vccd1 vccd1 _09020_ sky130_fd_sc_hd__xnor2_1
X_17389_ rbzero.debug_overlay.playerX\[3\] _01690_ _09620_ vssd1 vssd1 vccd1 vccd1
+ _01691_ sky130_fd_sc_hd__mux2_1
XFILLER_118_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18432__72 clknet_1_0__leaf__02438_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__inv_2
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10420_ rbzero.tex_b0\[57\] rbzero.tex_b0\[56\] _03269_ vssd1 vssd1 vccd1 vccd1 _03275_
+ sky130_fd_sc_hd__mux2_1
XFILLER_104_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10351_ rbzero.tex_b1\[25\] rbzero.tex_b1\[26\] _03232_ vssd1 vssd1 vccd1 vccd1 _03239_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13070_ _05826_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__inv_2
X_10282_ rbzero.tex_b1\[58\] rbzero.tex_b1\[59\] _03199_ vssd1 vssd1 vccd1 vccd1 _03203_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12021_ _04792_ net33 vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__nor2_1
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16760_ _09366_ _09367_ vssd1 vssd1 vccd1 vccd1 _09368_ sky130_fd_sc_hd__nor2_1
XFILLER_65_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13972_ _06719_ vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15711_ _08265_ _08392_ _08393_ vssd1 vssd1 vccd1 vccd1 _08394_ sky130_fd_sc_hd__o21ai_1
XFILLER_19_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12923_ _05678_ _05679_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__xnor2_1
X_16691_ _09298_ _09299_ vssd1 vssd1 vccd1 vccd1 _09300_ sky130_fd_sc_hd__xor2_1
XFILLER_46_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15642_ _07972_ _07959_ vssd1 vssd1 vccd1 vccd1 _08325_ sky130_fd_sc_hd__nor2_1
XFILLER_132_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _05609_ _05610_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__or2_1
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ net18 _04564_ _04576_ _04581_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__a31o_1
X_18361_ rbzero.pov.spi_counter\[5\] rbzero.pov.spi_counter\[4\] rbzero.pov.spi_counter\[3\]
+ rbzero.pov.spi_counter\[6\] vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__and4bb_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _08119_ _08122_ _08255_ vssd1 vssd1 vccd1 vccd1 _08257_ sky130_fd_sc_hd__nand3_1
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _05515_ _05534_ _05354_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__mux2_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17312_ _01628_ _01630_ _01629_ vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__o21ba_1
XFILLER_199_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14524_ _07193_ _07211_ vssd1 vssd1 vccd1 vccd1 _07212_ sky130_fd_sc_hd__xnor2_1
XFILLER_186_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18292_ _02378_ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__clkbuf_4
X_11736_ _04512_ _04513_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__and2_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17243_ _04986_ _01527_ _01577_ vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__a21oi_1
X_14455_ _07140_ _07142_ vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__xor2_1
XFILLER_186_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11667_ _03693_ _04445_ _04447_ _03669_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__o211a_1
XFILLER_179_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13406_ _06142_ _06154_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__xor2_1
XFILLER_127_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17174_ _01515_ _01516_ _01517_ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__and3_1
X_10618_ _03343_ _03390_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__xnor2_1
X_11598_ rbzero.tex_b0\[3\] rbzero.tex_b0\[2\] _04188_ vssd1 vssd1 vccd1 vccd1 _04380_
+ sky130_fd_sc_hd__mux2_1
X_14386_ _07064_ _07073_ vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__and2b_1
XFILLER_116_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16125_ _07265_ _08316_ vssd1 vssd1 vccd1 vccd1 _08738_ sky130_fd_sc_hd__and2_1
XFILLER_31_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13337_ _06090_ _06092_ _06093_ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__o21a_1
X_10549_ rbzero.map_rom.b6 vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__clkbuf_4
XFILLER_115_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16056_ _08668_ _08669_ vssd1 vssd1 vccd1 vccd1 _08670_ sky130_fd_sc_hd__and2_1
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13268_ _06023_ _06024_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__nor2_1
XFILLER_142_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15007_ _07571_ _07694_ _07573_ vssd1 vssd1 vccd1 vccd1 _07695_ sky130_fd_sc_hd__a21oi_1
X_12219_ rbzero.wall_tracer.trackDistX\[-7\] _04973_ _04974_ rbzero.wall_tracer.trackDistX\[-8\]
+ _04980_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__o221a_1
X_13199_ _05953_ _05955_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__or2_1
XFILLER_96_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19815_ clknet_leaf_2_i_clk _00746_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.ss_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16958_ _09443_ _09458_ _09456_ vssd1 vssd1 vccd1 vccd1 _09564_ sky130_fd_sc_hd__a21o_1
X_19746_ clknet_leaf_91_i_clk _00677_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15909_ rbzero.wall_tracer.trackDistX\[-9\] _08508_ _08525_ _08531_ vssd1 vssd1 vccd1
+ vccd1 _00540_ sky130_fd_sc_hd__o22a_1
X_19677_ clknet_leaf_81_i_clk _00608_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16889_ _09478_ _09479_ _09495_ vssd1 vssd1 vccd1 vccd1 _09496_ sky130_fd_sc_hd__a21o_1
XFILLER_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18628_ _02412_ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__clkbuf_4
XFILLER_64_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18559_ rbzero.pov.spi_buffer\[48\] rbzero.pov.spi_buffer\[49\] _02488_ vssd1 vssd1
+ vccd1 vccd1 _02498_ sky130_fd_sc_hd__mux2_1
XFILLER_75_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18922__107 clknet_1_0__leaf__02724_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__inv_2
XFILLER_33_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_12 _06899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 rbzero.spi_registers.vshift\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20521_ clknet_leaf_28_i_clk _01452_ vssd1 vssd1 vccd1 vccd1 gpout2.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_34 net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_45 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_56 _03338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_67 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20452_ net132 _01383_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20383_ net443 _01314_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12570_ _05310_ _05326_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__nand2_1
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11521_ _04301_ _04302_ _04303_ _03917_ _03689_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__o221a_1
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14240_ rbzero.debug_overlay.playerX\[-6\] _06888_ vssd1 vssd1 vccd1 vccd1 _06928_
+ sky130_fd_sc_hd__nand2_1
X_11452_ rbzero.color_sky\[3\] rbzero.color_floor\[3\] _03535_ vssd1 vssd1 vccd1 vccd1
+ _04235_ sky130_fd_sc_hd__mux2_1
XFILLER_109_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10403_ rbzero.tex_b1\[0\] rbzero.tex_b1\[1\] _02909_ vssd1 vssd1 vccd1 vccd1 _03266_
+ sky130_fd_sc_hd__mux2_1
XFILLER_171_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14171_ rbzero.wall_tracer.state\[13\] vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__inv_2
X_11383_ _04164_ _04165_ _04166_ _03740_ _03670_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__o221a_1
XFILLER_152_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10334_ rbzero.tex_b1\[33\] rbzero.tex_b1\[34\] _03221_ vssd1 vssd1 vccd1 vccd1 _03230_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13122_ _05433_ _05471_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__or2_1
XFILLER_194_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13053_ _05516_ _05496_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__nor2_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17930_ rbzero.pov.spi_buffer\[19\] rbzero.pov.ready_buffer\[19\] _02164_ vssd1 vssd1
+ vccd1 vccd1 _02165_ sky130_fd_sc_hd__mux2_1
X_10265_ rbzero.tex_g0\[3\] rbzero.tex_g0\[2\] _03188_ vssd1 vssd1 vccd1 vccd1 _03194_
+ sky130_fd_sc_hd__mux2_1
XFILLER_105_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12004_ net30 _04772_ _04775_ _04777_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__o211ai_1
XFILLER_3_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17861_ _02117_ _02119_ _02121_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__or3b_2
XFILLER_61_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10196_ rbzero.tex_g0\[36\] rbzero.tex_g0\[35\] _03155_ vssd1 vssd1 vccd1 vccd1 _03158_
+ sky130_fd_sc_hd__mux2_1
XFILLER_120_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19600_ clknet_leaf_26_i_clk _00531_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.wall\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_16812_ _09417_ _09418_ _09419_ vssd1 vssd1 vccd1 vccd1 _09420_ sky130_fd_sc_hd__or3_1
XFILLER_78_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17792_ _02056_ _02057_ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__nand2_1
XFILLER_4_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19531_ clknet_leaf_66_i_clk _00003_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16743_ _09264_ _09323_ _09350_ vssd1 vssd1 vccd1 vccd1 _09351_ sky130_fd_sc_hd__a21o_1
XFILLER_47_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13955_ _06637_ _06697_ _06698_ _06704_ vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__a31o_2
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12906_ _05661_ _05662_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__xnor2_1
X_19462_ clknet_leaf_56_i_clk _00408_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
X_16674_ _09282_ vssd1 vssd1 vccd1 vccd1 _09283_ sky130_fd_sc_hd__buf_2
XFILLER_34_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13886_ _06588_ _06572_ _06641_ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__a21o_1
XFILLER_59_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15625_ _08182_ _08308_ vssd1 vssd1 vccd1 vccd1 _08309_ sky130_fd_sc_hd__nor2_1
X_18411__53 clknet_1_1__leaf__02436_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__inv_2
X_12837_ _05499_ _05493_ _05593_ _05433_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__o22a_1
XFILLER_62_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19393_ rbzero.traced_texVinit\[0\] _08463_ _07815_ _08455_ vssd1 vssd1 vccd1 vccd1
+ _01428_ sky130_fd_sc_hd__a22o_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18344_ _02407_ vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__clkbuf_1
X_15556_ _08125_ _08223_ _08239_ vssd1 vssd1 vccd1 vccd1 _08240_ sky130_fd_sc_hd__a21o_1
XFILLER_15_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _05505_ _05470_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__nor2_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14507_ rbzero.wall_tracer.visualWallDist\[-10\] vssd1 vssd1 vccd1 vccd1 _07195_
+ sky130_fd_sc_hd__inv_2
X_18275_ rbzero.spi_registers.spi_cmd\[1\] _02981_ _02359_ _02107_ vssd1 vssd1 vccd1
+ vccd1 _02369_ sky130_fd_sc_hd__or4b_1
X_11719_ net8 _04495_ net4 _04496_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__and4b_1
XFILLER_175_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15487_ _08170_ _08171_ vssd1 vssd1 vccd1 vccd1 _08172_ sky130_fd_sc_hd__xor2_2
XFILLER_30_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12699_ _05394_ _05400_ _05274_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__mux2_1
X_17226_ _01560_ _01561_ _01562_ vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__or3_1
XFILLER_175_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14438_ _07124_ _07099_ vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__or2b_1
Xinput10 i_gpout1_sel[1] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_6
Xinput21 i_gpout3_sel[0] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__buf_4
Xinput32 i_gpout4_sel[5] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_4
XFILLER_122_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput43 i_reg_mosi vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_8
XFILLER_7_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17157_ _09675_ _01500_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14369_ _07005_ _07024_ _07037_ _07047_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__o22a_1
XFILLER_7_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16108_ _08719_ _08720_ vssd1 vssd1 vccd1 vccd1 _08721_ sky130_fd_sc_hd__nand2_2
XFILLER_116_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__02746_ clknet_0__02746_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02746_
+ sky130_fd_sc_hd__clkbuf_16
X_17088_ _09691_ _09692_ vssd1 vssd1 vccd1 vccd1 _09693_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16039_ _08651_ _08652_ vssd1 vssd1 vccd1 vccd1 _08653_ sky130_fd_sc_hd__nor2_1
XFILLER_69_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19729_ clknet_leaf_94_i_clk _00660_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19063__235 clknet_1_0__leaf__02737_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__inv_2
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20504_ clknet_leaf_42_i_clk _01435_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20435_ net495 _01366_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20366_ net426 _01297_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20297_ net357 _01228_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10050_ rbzero.tex_g1\[40\] rbzero.tex_g1\[41\] _03073_ vssd1 vssd1 vccd1 vccd1 _03081_
+ sky130_fd_sc_hd__mux2_1
XFILLER_121_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13740_ _06496_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__inv_2
X_10952_ _03736_ _03737_ _03677_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__mux2_1
XFILLER_43_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13671_ _06355_ _06380_ vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__nor2_1
X_10883_ _03634_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__buf_4
XFILLER_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15410_ _08002_ _07995_ vssd1 vssd1 vccd1 vccd1 _08095_ sky130_fd_sc_hd__or2b_1
XFILLER_31_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12622_ _05238_ _05349_ _05378_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__o21a_1
XFILLER_71_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16390_ _08985_ _09000_ vssd1 vssd1 vccd1 vccd1 _09001_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15341_ _08011_ _08025_ vssd1 vssd1 vccd1 vccd1 _08027_ sky130_fd_sc_hd__or2_1
XFILLER_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12553_ _05309_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__clkbuf_4
XFILLER_169_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11504_ _04285_ _04286_ _03917_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__mux2_1
XFILLER_129_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18060_ rbzero.spi_registers.spi_buffer\[6\] rbzero.spi_registers.spi_buffer\[5\]
+ _02227_ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__mux2_1
XFILLER_106_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15272_ _07956_ _07957_ vssd1 vssd1 vccd1 vccd1 _07958_ sky130_fd_sc_hd__nor2_1
X_12484_ _05119_ _05199_ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__nand2_1
XFILLER_184_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17011_ _09408_ vssd1 vssd1 vccd1 vccd1 _09617_ sky130_fd_sc_hd__inv_2
XFILLER_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14223_ rbzero.wall_tracer.visualWallDist\[-8\] _06910_ _03490_ vssd1 vssd1 vccd1
+ vccd1 _06911_ sky130_fd_sc_hd__mux2_1
X_11435_ rbzero.tex_g0\[43\] _03696_ _03697_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__and3_1
XFILLER_138_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14154_ _03485_ _06844_ vssd1 vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__and2_1
X_11366_ rbzero.color_sky\[2\] rbzero.color_floor\[2\] _03535_ vssd1 vssd1 vccd1 vccd1
+ _04150_ sky130_fd_sc_hd__mux2_1
XFILLER_153_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10317_ _03072_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__clkbuf_4
X_13105_ _05496_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__clkbuf_4
XFILLER_180_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_2_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11297_ _04035_ _04080_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__or2_2
X_14085_ rbzero.wall_tracer.visualWallDist\[3\] _06796_ _06785_ rbzero.wall_tracer.trackDistY\[3\]
+ _06797_ vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__o221a_1
XFILLER_152_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10248_ rbzero.tex_g0\[11\] rbzero.tex_g0\[10\] _03177_ vssd1 vssd1 vccd1 vccd1 _03185_
+ sky130_fd_sc_hd__mux2_1
X_13036_ _05789_ _05790_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__nor2_1
X_17913_ rbzero.pov.spi_buffer\[11\] rbzero.pov.ready_buffer\[11\] _02153_ vssd1 vssd1
+ vccd1 vccd1 _02156_ sky130_fd_sc_hd__mux2_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18893_ _02716_ vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17844_ rbzero.spi_registers.spi_counter\[1\] rbzero.spi_registers.spi_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__nand2_1
X_10179_ rbzero.tex_g0\[44\] rbzero.tex_g0\[43\] _03144_ vssd1 vssd1 vccd1 vccd1 _03149_
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17775_ _01985_ rbzero.debug_overlay.vplaneX\[-3\] vssd1 vssd1 vccd1 vccd1 _02042_
+ sky130_fd_sc_hd__nor2_1
X_14987_ _07668_ _07671_ _07674_ vssd1 vssd1 vccd1 vccd1 _07675_ sky130_fd_sc_hd__nor3_1
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16726_ _09332_ _09333_ vssd1 vssd1 vccd1 vccd1 _09334_ sky130_fd_sc_hd__xor2_1
X_19514_ clknet_leaf_52_i_clk _00460_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
X_13938_ _06603_ _06589_ _06653_ _05347_ vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__a211o_1
XFILLER_34_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19445_ gpout3.clk_div\[1\] gpout3.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__or2_1
X_16657_ _09264_ _09265_ vssd1 vssd1 vccd1 vccd1 _09266_ sky130_fd_sc_hd__nand2_1
X_13869_ _06619_ _06625_ _06603_ vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__mux2_1
X_15608_ _08289_ _08291_ vssd1 vssd1 vccd1 vccd1 _08292_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19376_ rbzero.traced_texa\[8\] rbzero.texV\[8\] vssd1 vssd1 vccd1 vccd1 _02854_
+ sky130_fd_sc_hd__or2_1
XFILLER_22_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16588_ rbzero.wall_tracer.trackDistX\[4\] rbzero.wall_tracer.stepDistX\[4\] vssd1
+ vssd1 vccd1 vccd1 _09198_ sky130_fd_sc_hd__nand2_1
XFILLER_15_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18327_ rbzero.spi_registers.new_other\[10\] rbzero.spi_registers.spi_buffer\[10\]
+ _02387_ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__mux2_1
XFILLER_176_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15539_ _08116_ _08127_ vssd1 vssd1 vccd1 vccd1 _08223_ sky130_fd_sc_hd__nand2_1
XFILLER_31_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18258_ rbzero.spi_registers.spi_done _02110_ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__nand2_1
XFILLER_147_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17209_ rbzero.wall_tracer.trackDistY\[-7\] rbzero.wall_tracer.stepDistY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__and2_1
XFILLER_191_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18189_ _04828_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__buf_2
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20220_ net280 _01151_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20151_ clknet_leaf_32_i_clk _01082_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[9\] sky130_fd_sc_hd__dfxtp_1
X_09962_ _03034_ vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__02729_ clknet_0__02729_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02729_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_131_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20082_ clknet_leaf_84_i_clk _01013_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
X_09893_ _02998_ vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__clkbuf_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18928__113 clknet_1_1__leaf__02724_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__inv_2
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11220_ _03886_ _03868_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__nand2_1
XFILLER_153_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20418_ net478 _01349_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18974__155 clknet_1_1__leaf__02728_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__inv_2
XFILLER_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11151_ _03733_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__buf_4
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20349_ net409 _01280_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10102_ _03108_ vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11082_ _03861_ _03863_ _03867_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__or3b_2
XFILLER_122_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10033_ _03071_ vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__clkbuf_1
X_14910_ _07594_ _07596_ _07597_ vssd1 vssd1 vccd1 vccd1 _07598_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15890_ _08512_ _08513_ _08514_ _08489_ vssd1 vssd1 vccd1 vccd1 _08515_ sky130_fd_sc_hd__a31o_1
XFILLER_102_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14841_ _07497_ _07522_ vssd1 vssd1 vccd1 vccd1 _07529_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17560_ _04109_ _01834_ vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__nand2_1
XFILLER_84_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14772_ _07447_ _07459_ vssd1 vssd1 vccd1 vccd1 _07460_ sky130_fd_sc_hd__xnor2_1
X_11984_ _04723_ _04749_ _04757_ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__a21boi_2
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16511_ _09111_ _09120_ vssd1 vssd1 vccd1 vccd1 _09121_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13723_ _05862_ _06156_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__nor2_1
X_10935_ _03624_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__buf_6
X_17491_ _01745_ _01775_ _01776_ _01783_ vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__a31o_1
XFILLER_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__02749_ clknet_0__02749_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02749_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_189_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16442_ _08807_ _09052_ vssd1 vssd1 vccd1 vccd1 _09053_ sky130_fd_sc_hd__xnor2_1
X_13654_ _06366_ _06410_ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10866_ _03610_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__buf_6
XFILLER_16_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12605_ _05258_ _05247_ _05313_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__mux2_1
X_16373_ _07972_ _08317_ vssd1 vssd1 vccd1 vccd1 _08984_ sky130_fd_sc_hd__and2_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13585_ _06336_ _06341_ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__or2b_1
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10797_ _03581_ _03577_ _03579_ vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__and3_1
XFILLER_13_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18112_ _03881_ _02263_ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__nand2_1
X_15324_ _08008_ _08009_ vssd1 vssd1 vccd1 vccd1 _08010_ sky130_fd_sc_hd__and2_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12536_ _05252_ _05287_ _05292_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__and3_1
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18043_ _02223_ vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__clkbuf_1
X_15255_ _07782_ _07792_ _07849_ _07847_ vssd1 vssd1 vccd1 vccd1 _07941_ sky130_fd_sc_hd__a31o_2
X_12467_ _05158_ _05221_ _05222_ _05223_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__or4_4
XFILLER_172_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14206_ _03490_ rbzero.wall_tracer.stepDistY\[-4\] _04947_ vssd1 vssd1 vccd1 vccd1
+ _06894_ sky130_fd_sc_hd__a21oi_1
X_11418_ rbzero.tex_g0\[61\] rbzero.tex_g0\[60\] _03700_ vssd1 vssd1 vccd1 vccd1 _04202_
+ sky130_fd_sc_hd__mux2_1
XFILLER_193_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15186_ _07871_ _07872_ vssd1 vssd1 vccd1 vccd1 _07873_ sky130_fd_sc_hd__nand2_1
X_12398_ _03488_ _05078_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__or2_1
X_19092__261 clknet_1_0__leaf__02740_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__inv_2
XFILLER_99_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14137_ _06833_ vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__clkbuf_1
XFILLER_153_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11349_ rbzero.debug_overlay.playerX\[-2\] _04056_ _04128_ _04133_ vssd1 vssd1 vccd1
+ vccd1 _04134_ sky130_fd_sc_hd__a211o_1
X_19994_ clknet_leaf_94_i_clk _00925_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14068_ _03484_ vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__clkbuf_4
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13019_ _05775_ _05743_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__xnor2_1
XFILLER_95_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18876_ _04500_ _02286_ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__nand2_1
XFILLER_67_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17827_ _02088_ _02089_ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__nand2_1
XFILLER_66_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17758_ _01972_ _04102_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__xor2_1
XFILLER_130_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16709_ _09220_ _09221_ _09224_ vssd1 vssd1 vccd1 vccd1 _09317_ sky130_fd_sc_hd__o21ba_1
X_17689_ rbzero.debug_overlay.vplaneX\[-1\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__nand2_1
XFILLER_74_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19428_ _01925_ _02883_ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19359_ rbzero.traced_texa\[5\] rbzero.texV\[5\] vssd1 vssd1 vccd1 vccd1 _02840_
+ sky130_fd_sc_hd__nor2_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19175__336 clknet_1_1__leaf__02748_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__inv_2
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20203_ net263 _01134_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20134_ clknet_leaf_89_i_clk _01065_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_104_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09945_ _03025_ vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18439__78 clknet_1_1__leaf__02439_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__inv_2
XFILLER_132_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20065_ clknet_leaf_83_i_clk _00996_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_58_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09876_ _02989_ vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__clkbuf_1
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10720_ _03484_ _03507_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__and2_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10651_ rbzero.map_overlay.i_mapdy\[3\] vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__inv_2
XFILLER_201_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13370_ _06097_ _06121_ _06056_ _06126_ vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__o31a_1
X_10582_ rbzero.debug_overlay.playerX\[5\] vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__inv_2
XFILLER_155_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12321_ _04877_ _04878_ _04879_ _04880_ _03479_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__o311a_4
XFILLER_5_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15040_ _07096_ _07098_ _07095_ vssd1 vssd1 vccd1 vccd1 _07728_ sky130_fd_sc_hd__a21bo_1
XFILLER_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12252_ _05007_ _05011_ _05012_ _05009_ rbzero.wall_tracer.mapY\[7\] vssd1 vssd1
+ vccd1 vccd1 _00402_ sky130_fd_sc_hd__a32o_1
XFILLER_107_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11203_ rbzero.tex_r1\[21\] _03660_ _03768_ _03702_ vssd1 vssd1 vccd1 vccd1 _03988_
+ sky130_fd_sc_hd__a31o_1
X_12183_ _04926_ _04930_ _04944_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__or3_1
XFILLER_107_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11134_ _03823_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__clkbuf_4
X_16991_ _09595_ _09596_ vssd1 vssd1 vccd1 vccd1 _09597_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_82_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_110_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18730_ _02610_ _02611_ vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__nand2_1
XFILLER_62_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11065_ gpout0.vpos\[6\] _03447_ rbzero.map_overlay.i_mapdy\[2\] _03849_ _03850_
+ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__o221a_1
X_15942_ rbzero.wall_tracer.trackDistX\[-5\] _08553_ _08554_ _08560_ vssd1 vssd1 vccd1
+ vccd1 _00544_ sky130_fd_sc_hd__o22a_1
XFILLER_27_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10016_ rbzero.tex_g1\[56\] rbzero.tex_g1\[57\] _03061_ vssd1 vssd1 vccd1 vccd1 _03063_
+ sky130_fd_sc_hd__mux2_1
X_18661_ rbzero.debug_overlay.playerX\[-1\] _02534_ _02558_ _02559_ vssd1 vssd1 vccd1
+ vccd1 _01004_ sky130_fd_sc_hd__a211o_1
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ _08498_ _08499_ vssd1 vssd1 vccd1 vccd1 _08500_ sky130_fd_sc_hd__xnor2_1
XFILLER_92_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17612_ _01894_ _03390_ _05009_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__mux2_1
XFILLER_91_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14824_ _07502_ _07510_ _07511_ vssd1 vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__a21o_1
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18592_ _02515_ vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__clkbuf_1
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17543_ _01829_ _01830_ _01831_ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__nand3_1
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14755_ _07433_ _07440_ _07442_ vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__a21oi_2
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ _04736_ _04739_ _04740_ net32 vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__or4b_1
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13706_ _06451_ _06462_ vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__xor2_1
X_10918_ _03627_ vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__buf_4
X_17474_ _01765_ _01766_ _01764_ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__a21o_1
XFILLER_189_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_14686_ _07373_ _07360_ vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__xnor2_1
X_11898_ _03459_ _03469_ _04672_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__mux2_1
X_16425_ _08391_ vssd1 vssd1 vccd1 vccd1 _09036_ sky130_fd_sc_hd__clkbuf_4
XFILLER_34_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13637_ _06389_ _06393_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__xnor2_1
X_10849_ _03558_ _03603_ _03608_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__nor3b_4
XFILLER_13_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16356_ _08725_ _08950_ _08949_ vssd1 vssd1 vccd1 vccd1 _08967_ sky130_fd_sc_hd__a21o_1
XFILLER_158_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13568_ _06308_ _06323_ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__nor2_1
XFILLER_185_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15307_ _07123_ vssd1 vssd1 vccd1 vccd1 _07993_ sky130_fd_sc_hd__clkbuf_4
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12519_ _05234_ _05238_ _05275_ _05246_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__o31a_2
XFILLER_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16287_ _08252_ vssd1 vssd1 vccd1 vccd1 _08899_ sky130_fd_sc_hd__buf_2
XFILLER_145_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_35_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13499_ _06174_ _06170_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__and2b_1
XFILLER_173_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18026_ rbzero.pov.spi_buffer\[65\] rbzero.pov.ready_buffer\[65\] _02208_ vssd1 vssd1
+ vccd1 vccd1 _02215_ sky130_fd_sc_hd__mux2_1
XFILLER_117_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15238_ _07799_ _07801_ vssd1 vssd1 vccd1 vccd1 _07925_ sky130_fd_sc_hd__nor2_1
XFILLER_160_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15169_ _07007_ vssd1 vssd1 vccd1 vccd1 _07856_ sky130_fd_sc_hd__buf_2
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19977_ net206 _00908_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09730_ _02911_ vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18859_ _02415_ _02414_ _02420_ rbzero.pov.spi_done vssd1 vssd1 vccd1 vccd1 _02692_
+ sky130_fd_sc_hd__a31o_1
XFILLER_95_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19099__267 clknet_1_1__leaf__02741_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__inv_2
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20117_ clknet_leaf_76_i_clk _01048_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_104_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09928_ _03016_ vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20048_ clknet_leaf_81_i_clk _00979_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[64\]
+ sky130_fd_sc_hd__dfxtp_1
X_09859_ rbzero.tex_r1\[1\] rbzero.tex_r1\[2\] _02976_ vssd1 vssd1 vccd1 vccd1 _02979_
+ sky130_fd_sc_hd__mux2_1
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _05614_ _05626_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ net50 _04566_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__and2_1
XFILLER_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _07219_ _07226_ _07227_ vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__a21boi_1
XFILLER_183_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _03537_ _04515_ _04516_ net40 _04529_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__a221o_1
XFILLER_198_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _03491_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__buf_4
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ rbzero.wall_tracer.stepDistY\[3\] vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__inv_2
X_11683_ rbzero.tex_b1\[2\] _03690_ _03823_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__a21o_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16210_ _08821_ _08822_ vssd1 vssd1 vccd1 vccd1 _08823_ sky130_fd_sc_hd__nor2_1
X_13422_ _06176_ _06178_ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__and2_1
X_10634_ rbzero.map_overlay.i_otherx\[1\] vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__inv_2
X_17190_ _01529_ _01530_ _01524_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__a21bo_1
XFILLER_201_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19158__320 clknet_1_0__leaf__02747_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__inv_2
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16141_ _08752_ _08753_ vssd1 vssd1 vccd1 vccd1 _08754_ sky130_fd_sc_hd__nand2_1
XFILLER_128_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13353_ _05609_ _06011_ _06015_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__and3b_1
X_10565_ rbzero.debug_overlay.playerY\[4\] _03359_ rbzero.wall_tracer.mapY\[5\] _03360_
+ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__a22o_1
XFILLER_6_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12304_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[10\] vssd1
+ vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__nor2_1
X_16072_ _08679_ _08685_ vssd1 vssd1 vccd1 vccd1 _08686_ sky130_fd_sc_hd__xor2_1
X_13284_ _05609_ _06016_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__or2_1
X_10496_ rbzero.tex_b0\[21\] rbzero.tex_b0\[20\] _03313_ vssd1 vssd1 vccd1 vccd1 _03315_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15023_ _07265_ _07270_ vssd1 vssd1 vccd1 vccd1 _07711_ sky130_fd_sc_hd__nor2_1
X_19900_ clknet_leaf_16_i_clk _00831_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_136_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12235_ _04960_ rbzero.wall_tracer.trackDistX\[4\] _04961_ rbzero.wall_tracer.trackDistX\[3\]
+ _04996_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__a221o_1
XFILLER_64_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19831_ clknet_leaf_4_i_clk _00762_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12166_ _04927_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__clkbuf_4
XFILLER_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11117_ _03902_ _03834_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__nand2_1
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19762_ clknet_leaf_86_i_clk _00693_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_16974_ _09579_ _09483_ _09480_ vssd1 vssd1 vccd1 vccd1 _09580_ sky130_fd_sc_hd__a21o_1
X_18418__59 clknet_1_1__leaf__02437_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__inv_2
X_12097_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__nand2_1
XFILLER_111_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18713_ rbzero.pov.ready_buffer\[49\] _02413_ _02582_ _02599_ vssd1 vssd1 vccd1 vccd1
+ _02600_ sky130_fd_sc_hd__a211o_1
XFILLER_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11048_ gpout0.vpos\[4\] vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__buf_4
X_15925_ rbzero.wall_tracer.trackDistX\[-7\] _08508_ _08539_ _08545_ vssd1 vssd1 vccd1
+ vccd1 _00542_ sky130_fd_sc_hd__o22a_1
X_19693_ clknet_leaf_9_i_clk _00624_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.i_row\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_76_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput8 i_gpout0_sel[5] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_6
XFILLER_49_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18644_ rbzero.debug_overlay.playerX\[-6\] _02542_ vssd1 vssd1 vccd1 vccd1 _02548_
+ sky130_fd_sc_hd__or2_1
X_15856_ _04951_ _04952_ _06784_ vssd1 vssd1 vccd1 vccd1 _08486_ sky130_fd_sc_hd__or3b_1
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14807_ _06872_ _07494_ _07273_ _06866_ vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__o22a_1
XFILLER_188_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18575_ _02506_ vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__clkbuf_1
X_15787_ _08452_ vssd1 vssd1 vccd1 vccd1 _08455_ sky130_fd_sc_hd__buf_2
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12999_ _05718_ _05720_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__xor2_1
XFILLER_45_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17526_ _01814_ _01801_ _01815_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__a21oi_1
X_14738_ _07415_ _07420_ _07419_ vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__o21ba_1
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17457_ rbzero.debug_overlay.vplaneY\[-9\] vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__inv_2
X_14669_ _07342_ _07354_ vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__nor2_1
X_16408_ _08108_ _08130_ vssd1 vssd1 vccd1 vccd1 _09019_ sky130_fd_sc_hd__or2_1
X_17388_ _08478_ _01689_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__xnor2_1
XFILLER_192_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16339_ _08949_ _08950_ vssd1 vssd1 vccd1 vccd1 _08951_ sky130_fd_sc_hd__and2b_1
XFILLER_146_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18009_ rbzero.pov.spi_buffer\[57\] rbzero.pov.ready_buffer\[57\] _02197_ vssd1 vssd1
+ vccd1 vccd1 _02206_ sky130_fd_sc_hd__mux2_1
XFILLER_161_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10350_ _03238_ vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10281_ _03202_ vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12020_ net44 _04792_ _04790_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__and3_1
XFILLER_183_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13971_ rbzero.wall_tracer.stepDistY\[-2\] _06717_ _06718_ vssd1 vssd1 vccd1 vccd1
+ _06719_ sky130_fd_sc_hd__mux2_1
X_15710_ _07662_ _08018_ _08391_ _07213_ vssd1 vssd1 vccd1 vccd1 _08393_ sky130_fd_sc_hd__o22ai_1
XFILLER_58_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12922_ _05571_ _05572_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__xnor2_1
X_16690_ _09097_ _09184_ _09183_ vssd1 vssd1 vccd1 vccd1 _09299_ sky130_fd_sc_hd__a21oi_1
XFILLER_150_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15641_ _08242_ _08222_ vssd1 vssd1 vccd1 vccd1 _08324_ sky130_fd_sc_hd__or2b_1
XFILLER_62_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12853_ _05546_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__clkbuf_4
XFILLER_34_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ net44 _04568_ _04577_ _04578_ _04580_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__a311o_1
X_18360_ rbzero.pov.spi_counter\[0\] _02414_ rbzero.pov.spi_counter\[1\] vssd1 vssd1
+ vccd1 vccd1 _02418_ sky130_fd_sc_hd__a21o_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15572_ _08119_ _08122_ _08255_ vssd1 vssd1 vccd1 vccd1 _08256_ sky130_fd_sc_hd__a21o_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _05392_ _05536_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__nor2_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _01634_ _01635_ vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__and2b_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _07154_ _07178_ _07200_ _07196_ _07194_ vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__o32a_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18291_ _02107_ _01658_ _02981_ _02359_ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__or4_1
X_11735_ net6 _04496_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__nor2_2
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _08485_ _01575_ _01576_ _08575_ _01522_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__o311a_1
X_14454_ _07100_ _07141_ vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__nor2_1
XFILLER_41_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11666_ _03823_ _04446_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__or2_1
XFILLER_174_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13405_ _06158_ _06161_ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__or2_1
X_17173_ rbzero.wall_tracer.trackDistX\[10\] rbzero.wall_tracer.stepDistX\[10\] vssd1
+ vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__nand2_1
X_10617_ _03369_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__inv_2
X_14385_ _07065_ _07069_ _07072_ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__o21ai_1
XFILLER_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11597_ rbzero.tex_b0\[1\] rbzero.tex_b0\[0\] _04188_ vssd1 vssd1 vccd1 vccd1 _04379_
+ sky130_fd_sc_hd__mux2_1
X_16124_ _08735_ _08736_ vssd1 vssd1 vccd1 vccd1 _08737_ sky130_fd_sc_hd__xor2_1
X_13336_ _06058_ _06089_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__nand2_1
XFILLER_116_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10548_ rbzero.debug_overlay.playerY\[4\] vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__inv_2
XFILLER_143_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16055_ _08662_ _08667_ vssd1 vssd1 vccd1 vccd1 _08669_ sky130_fd_sc_hd__or2_1
XFILLER_157_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13267_ _05957_ _06006_ _06022_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__nor3_1
X_10479_ rbzero.tex_b0\[29\] rbzero.tex_b0\[28\] _03302_ vssd1 vssd1 vccd1 vccd1 _03306_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15006_ _07572_ _07610_ vssd1 vssd1 vccd1 vccd1 _07694_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12218_ _04974_ rbzero.wall_tracer.trackDistX\[-8\] _04975_ rbzero.wall_tracer.trackDistX\[-9\]
+ _04979_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__a221o_1
XFILLER_194_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13198_ _05480_ _05954_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__nor2_1
XFILLER_123_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19814_ clknet_leaf_1_i_clk _00745_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.ss_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12149_ _04909_ _04910_ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__nand2_1
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19745_ clknet_leaf_91_i_clk _00676_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16957_ _09561_ _09562_ vssd1 vssd1 vccd1 vccd1 _09563_ sky130_fd_sc_hd__xor2_1
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15908_ _08512_ _08529_ _08530_ _08522_ vssd1 vssd1 vccd1 vccd1 _08531_ sky130_fd_sc_hd__a31o_1
X_19676_ clknet_leaf_79_i_clk _00607_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
X_16888_ _09493_ _09494_ vssd1 vssd1 vccd1 vccd1 _09495_ sky130_fd_sc_hd__nand2_1
XFILLER_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18627_ _02533_ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__clkbuf_4
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15839_ _03364_ _07936_ vssd1 vssd1 vccd1 vccd1 _08469_ sky130_fd_sc_hd__nor2_1
XFILLER_80_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18558_ _02497_ vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17509_ _01784_ rbzero.wall_tracer.rayAddendY\[3\] vssd1 vssd1 vccd1 vccd1 _01800_
+ sky130_fd_sc_hd__nor2_1
XFILLER_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18489_ _02461_ vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_13 _06938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20520_ clknet_leaf_42_i_clk _01451_ vssd1 vssd1 vccd1 vccd1 gpout2.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_24 rbzero.wall_tracer.rayAddendX\[-3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_35 net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_46 net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_57 _03688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20451_ net131 _01382_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[42\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_68 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20382_ net442 _01313_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_180_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19040__214 clknet_1_0__leaf__02735_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__inv_2
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11520_ rbzero.tex_g1\[45\] rbzero.tex_g1\[44\] _03727_ vssd1 vssd1 vccd1 vccd1 _04303_
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11451_ _04234_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__buf_4
X_10402_ _03265_ vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14170_ _06857_ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__buf_2
X_11382_ rbzero.tex_g0\[29\] rbzero.tex_g0\[28\] _03709_ vssd1 vssd1 vccd1 vccd1 _04166_
+ sky130_fd_sc_hd__mux2_1
XFILLER_165_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13121_ _05484_ _05517_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__or2_1
X_10333_ _03229_ vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13052_ _05804_ _05808_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__nand2_1
X_10264_ _03193_ vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12003_ _04750_ net67 _04776_ net31 vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__a211o_1
XFILLER_121_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10195_ _03157_ vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__clkbuf_1
X_17860_ rbzero.spi_registers.spi_counter\[3\] rbzero.spi_registers.spi_counter\[0\]
+ _02120_ _02109_ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__a31o_1
XFILLER_132_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16811_ _09309_ _09311_ _09310_ vssd1 vssd1 vccd1 vccd1 _09419_ sky130_fd_sc_hd__o21ba_1
X_17791_ rbzero.debug_overlay.vplaneX\[-2\] _02042_ vssd1 vssd1 vccd1 vccd1 _02057_
+ sky130_fd_sc_hd__nand2_1
X_19530_ clknet_leaf_62_i_clk _00002_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16742_ _09348_ _09349_ vssd1 vssd1 vccd1 vccd1 _09350_ sky130_fd_sc_hd__nand2_1
XFILLER_19_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13954_ _05476_ _06703_ _06629_ vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__a21o_1
XFILLER_98_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12905_ _05525_ _05518_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__xnor2_1
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16673_ _09280_ _09281_ vssd1 vssd1 vccd1 vccd1 _09282_ sky130_fd_sc_hd__and2_1
XFILLER_62_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19461_ clknet_leaf_54_i_clk _00407_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13885_ _06588_ _06620_ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__nor2_1
XFILLER_28_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12836_ _05592_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__buf_2
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15624_ _07937_ _08307_ vssd1 vssd1 vccd1 vccd1 _08308_ sky130_fd_sc_hd__xnor2_1
X_19392_ rbzero.texV\[10\] _02762_ _02709_ _02867_ vssd1 vssd1 vccd1 vccd1 _01427_
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15555_ _08228_ _08238_ vssd1 vssd1 vccd1 vccd1 _08239_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18343_ rbzero.spi_registers.new_vshift\[5\] rbzero.spi_registers.spi_buffer\[5\]
+ _02401_ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__mux2_1
X_12767_ _05501_ _05512_ _05523_ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__o21a_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _06787_ _04840_ _06860_ _07152_ vssd1 vssd1 vccd1 vccd1 _07194_ sky130_fd_sc_hd__and4_1
X_18274_ rbzero.spi_registers.got_new_sky _02285_ _02283_ _02368_ vssd1 vssd1 vccd1
+ vccd1 _00808_ sky130_fd_sc_hd__a31o_1
X_11718_ net5 vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__buf_2
XFILLER_175_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15486_ _07941_ _08044_ _08042_ vssd1 vssd1 vccd1 vccd1 _08171_ sky130_fd_sc_hd__a21oi_2
XFILLER_159_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12698_ _05357_ _05395_ _05410_ _05365_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__a22o_1
XFILLER_147_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14437_ _07099_ _07124_ vssd1 vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__or2b_1
X_17225_ _01553_ _01555_ _01554_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__a21boi_1
X_11649_ _03693_ _04427_ _04429_ _03669_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__o211a_1
Xinput11 i_gpout1_sel[2] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_6
XFILLER_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 i_gpout3_sel[1] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_4
Xinput33 i_gpout5_sel[0] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__buf_4
X_17156_ _08889_ _09035_ vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__nor2_1
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput44 i_reg_sclk vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__buf_8
X_14368_ _07024_ _07038_ _07047_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__nor3_1
XFILLER_183_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16107_ _08598_ _08709_ vssd1 vssd1 vccd1 vccd1 _08720_ sky130_fd_sc_hd__nand2_1
XFILLER_116_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13319_ _06073_ _06075_ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__nor2_1
X_17087_ _09561_ _09562_ _09599_ vssd1 vssd1 vccd1 vccd1 _09692_ sky130_fd_sc_hd__o21a_1
Xclkbuf_1_1__f__02745_ clknet_0__02745_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02745_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_182_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14299_ rbzero.debug_overlay.playerX\[-3\] _06961_ vssd1 vssd1 vccd1 vccd1 _06987_
+ sky130_fd_sc_hd__or2_1
XFILLER_115_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16038_ _08365_ _08368_ _08367_ vssd1 vssd1 vccd1 vccd1 _08652_ sky130_fd_sc_hd__a21boi_1
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17989_ _02195_ vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19728_ clknet_leaf_94_i_clk _00659_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19659_ clknet_leaf_15_i_clk _00590_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20503_ clknet_leaf_42_i_clk _01434_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_194_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20434_ net494 _01365_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20365_ net425 _01296_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20296_ net356 _01227_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10951_ rbzero.tex_r0\[35\] rbzero.tex_r0\[34\] _03663_ vssd1 vssd1 vccd1 vccd1 _03737_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13670_ _06304_ _06327_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__xnor2_1
XFILLER_189_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10882_ _03666_ _03667_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__or2_1
X_12621_ _05244_ _05276_ _05297_ _05212_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__a31o_1
XFILLER_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15340_ _08011_ _08025_ vssd1 vssd1 vccd1 vccd1 _08026_ sky130_fd_sc_hd__nand2_1
XFILLER_24_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12552_ _05300_ _05308_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__nand2_1
XFILLER_185_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11503_ rbzero.tex_g1\[59\] rbzero.tex_g1\[58\] _03727_ vssd1 vssd1 vccd1 vccd1 _04286_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15271_ _07953_ _07955_ vssd1 vssd1 vccd1 vccd1 _07957_ sky130_fd_sc_hd__and2_1
XFILLER_12_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12483_ _05118_ _05239_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__xnor2_1
X_17010_ _09092_ _09411_ _09412_ vssd1 vssd1 vccd1 vccd1 _09616_ sky130_fd_sc_hd__a21o_1
XFILLER_156_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14222_ rbzero.debug_overlay.playerY\[-8\] _06909_ _04928_ vssd1 vssd1 vccd1 vccd1
+ _06910_ sky130_fd_sc_hd__mux2_1
X_11434_ rbzero.tex_g0\[41\] rbzero.tex_g0\[40\] _04188_ vssd1 vssd1 vccd1 vccd1 _04218_
+ sky130_fd_sc_hd__mux2_1
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14153_ _06843_ rbzero.wall_tracer.wall\[0\] _03458_ vssd1 vssd1 vccd1 vccd1 _06844_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11365_ _04149_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__buf_4
XFILLER_180_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13104_ _05301_ _05610_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__nor2_1
X_10316_ _03220_ vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14084_ rbzero.wall_tracer.trackDistX\[2\] _06788_ _06805_ vssd1 vssd1 vccd1 vccd1
+ _00441_ sky130_fd_sc_hd__o21a_1
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11296_ _04074_ _04080_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__nor2_4
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _05770_ _05773_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__or2b_1
X_17912_ _02155_ vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__clkbuf_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10247_ _03184_ vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18892_ _02714_ _04834_ _02715_ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__and3b_1
X_18951__134 clknet_1_1__leaf__02726_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__inv_2
XFILLER_152_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17843_ rbzero.spi_registers.spi_counter\[0\] vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__inv_2
XFILLER_113_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10178_ _03148_ vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17774_ _02039_ _02037_ _02038_ _08464_ vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__a31o_1
X_14986_ _07655_ _07669_ _07672_ _07673_ vssd1 vssd1 vccd1 vccd1 _07674_ sky130_fd_sc_hd__o211a_1
X_19513_ clknet_leaf_53_i_clk _00459_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16725_ _08107_ _08317_ vssd1 vssd1 vccd1 vccd1 _09333_ sky130_fd_sc_hd__and2_1
XFILLER_47_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13937_ _05325_ _06602_ _06651_ _05271_ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__a211o_1
XFILLER_62_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19444_ gpout3.clk_div\[1\] gpout3.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__nand2_1
X_16656_ _09161_ _09247_ _09263_ vssd1 vssd1 vccd1 vccd1 _09265_ sky130_fd_sc_hd__nand3_1
X_13868_ _06621_ _06624_ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__nor2_1
XFILLER_50_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15607_ _08093_ _08165_ _08290_ vssd1 vssd1 vccd1 vccd1 _08291_ sky130_fd_sc_hd__a21oi_1
X_12819_ _05450_ _05545_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__nand2_2
XFILLER_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19375_ rbzero.texV\[7\] _02762_ _02709_ _02853_ vssd1 vssd1 vccd1 vccd1 _01424_
+ sky130_fd_sc_hd__a22o_1
X_16587_ _08485_ _09195_ _09196_ vssd1 vssd1 vccd1 vccd1 _09197_ sky130_fd_sc_hd__and3_2
X_13799_ _06477_ _06508_ _06511_ _06543_ _06555_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__o221a_1
XFILLER_16_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18326_ _02397_ vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__clkbuf_1
X_15538_ _08101_ _08112_ _08110_ vssd1 vssd1 vccd1 vccd1 _08222_ sky130_fd_sc_hd__a21o_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15469_ _08129_ _08026_ _08153_ vssd1 vssd1 vccd1 vccd1 _08154_ sky130_fd_sc_hd__a21oi_1
X_18257_ _02358_ vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17208_ rbzero.wall_tracer.trackDistY\[-7\] rbzero.wall_tracer.stepDistY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__nor2_1
XFILLER_163_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18188_ rbzero.floor_leak\[1\] _02311_ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__or2_1
XFILLER_162_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17139_ _09009_ _09046_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__nor2_1
XFILLER_143_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20150_ clknet_leaf_20_i_clk _01081_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[8\] sky130_fd_sc_hd__dfxtp_1
X_09961_ rbzero.tex_r0\[19\] rbzero.tex_r0\[18\] _03028_ vssd1 vssd1 vccd1 vccd1 _03034_
+ sky130_fd_sc_hd__mux2_1
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__02728_ clknet_0__02728_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02728_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_171_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20081_ clknet_leaf_84_i_clk _01012_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
X_09892_ rbzero.tex_r0\[52\] rbzero.tex_r0\[51\] _02995_ vssd1 vssd1 vccd1 vccd1 _02998_
+ sky130_fd_sc_hd__mux2_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18387__31 clknet_1_0__leaf__02434_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__inv_2
XFILLER_20_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20417_ net477 _01348_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19152__315 clknet_1_0__leaf__02746_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__inv_2
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11150_ rbzero.tex_r1\[59\] _03925_ _03934_ _03726_ vssd1 vssd1 vccd1 vccd1 _03935_
+ sky130_fd_sc_hd__o211a_1
XFILLER_190_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20348_ net408 _01279_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[3\] sky130_fd_sc_hd__dfxtp_1
X_10101_ rbzero.tex_g1\[16\] rbzero.tex_g1\[17\] _03106_ vssd1 vssd1 vccd1 vccd1 _03108_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11081_ _03425_ _03523_ _02900_ _03864_ _03866_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__o221a_1
X_20279_ net339 _01210_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10032_ rbzero.tex_g1\[48\] rbzero.tex_g1\[49\] _03061_ vssd1 vssd1 vccd1 vccd1 _03071_
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14840_ _07477_ _07527_ vssd1 vssd1 vccd1 vccd1 _07528_ sky130_fd_sc_hd__xnor2_2
XFILLER_29_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14771_ _07448_ _07454_ _07458_ vssd1 vssd1 vccd1 vccd1 _07459_ sky130_fd_sc_hd__o21ai_1
X_11983_ net28 _04752_ _04754_ _04756_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__a31o_1
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16510_ _09118_ _09119_ vssd1 vssd1 vccd1 vccd1 _09120_ sky130_fd_sc_hd__nor2_1
X_13722_ _06443_ _06459_ _06460_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__a21o_1
X_10934_ _03688_ _03705_ _03714_ _03719_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__a31o_1
XFILLER_17_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17490_ rbzero.wall_tracer.rayAddendY\[1\] _08447_ _01782_ _01714_ vssd1 vssd1 vccd1
+ vccd1 _01783_ sky130_fd_sc_hd__a22o_1
XFILLER_90_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__02748_ clknet_0__02748_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02748_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16441_ _09046_ _09050_ _09051_ vssd1 vssd1 vccd1 vccd1 _09052_ sky130_fd_sc_hd__o21a_1
X_13653_ _06121_ _05994_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__nor2_1
X_10865_ rbzero.tex_r0\[5\] rbzero.tex_r0\[4\] _03649_ vssd1 vssd1 vccd1 vccd1 _03651_
+ sky130_fd_sc_hd__mux2_1
XFILLER_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12604_ _05360_ _05225_ _05311_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__mux2_1
X_16372_ _08981_ _08982_ vssd1 vssd1 vccd1 vccd1 _08983_ sky130_fd_sc_hd__nor2_1
XFILLER_176_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13584_ _06125_ _06337_ _06339_ _06340_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__a22o_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ _03577_ _03579_ _03581_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__a21oi_1
XFILLER_157_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15323_ _07617_ _07748_ _07756_ _07646_ vssd1 vssd1 vccd1 vccd1 _08009_ sky130_fd_sc_hd__o22ai_1
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18111_ _02263_ vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__buf_2
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12535_ _05198_ _05201_ _05291_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__o21ai_1
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15254_ _07924_ _07926_ vssd1 vssd1 vccd1 vccd1 _07940_ sky130_fd_sc_hd__nor2_2
XFILLER_8_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18042_ rbzero.pov.spi_buffer\[73\] rbzero.pov.ready_buffer\[73\] _02142_ vssd1 vssd1
+ vccd1 vccd1 _02223_ sky130_fd_sc_hd__mux2_1
XFILLER_173_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12466_ _05161_ _05183_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__xnor2_2
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14205_ _04947_ _06881_ _06891_ _06892_ vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__a2bb2o_4
X_11417_ _04199_ _04200_ _03740_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__mux2_1
X_15185_ _07738_ _07852_ _07870_ vssd1 vssd1 vccd1 vccd1 _07872_ sky130_fd_sc_hd__nand3_1
XFILLER_153_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12397_ _05077_ _05150_ _05153_ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__a21oi_1
XFILLER_126_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14136_ rbzero.wall_tracer.stepDistX\[5\] _06765_ _06825_ vssd1 vssd1 vccd1 vccd1
+ _06833_ sky130_fd_sc_hd__mux2_1
XFILLER_152_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11348_ rbzero.debug_overlay.playerX\[1\] _04066_ _04129_ _04132_ vssd1 vssd1 vccd1
+ vccd1 _04133_ sky130_fd_sc_hd__a211o_1
XFILLER_180_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19993_ clknet_leaf_95_i_clk _00924_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14067_ _03495_ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__clkbuf_4
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11279_ _04051_ _04063_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__nor2_1
X_13018_ _05744_ _05740_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__and2b_1
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18875_ _02704_ vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17826_ _02001_ rbzero.wall_tracer.rayAddendX\[9\] vssd1 vssd1 vccd1 vccd1 _02089_
+ sky130_fd_sc_hd__nand2_1
XFILLER_39_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17757_ _08458_ _02014_ _02015_ _02025_ vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__a31o_1
XFILLER_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14969_ _07006_ _07157_ _07178_ _07048_ vssd1 vssd1 vccd1 vccd1 _07657_ sky130_fd_sc_hd__o22a_1
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16708_ _09244_ _09211_ vssd1 vssd1 vccd1 vccd1 _09316_ sky130_fd_sc_hd__or2b_1
X_17688_ rbzero.debug_overlay.vplaneX\[-1\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__or2_1
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19427_ _01920_ _01926_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__and2b_1
XFILLER_35_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16639_ _06858_ _07012_ _08130_ _09142_ vssd1 vssd1 vccd1 vccd1 _09248_ sky130_fd_sc_hd__or4_1
XFILLER_50_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19358_ _02834_ _02836_ _02835_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__a21boi_1
XFILLER_149_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18309_ rbzero.spi_registers.new_other\[0\] rbzero.spi_registers.spi_buffer\[0\]
+ _02388_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__mux2_1
XFILLER_200_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19289_ _02759_ _02780_ _02781_ _02762_ rbzero.texV\[-7\] vssd1 vssd1 vccd1 vccd1
+ _01410_ sky130_fd_sc_hd__a32o_1
X_19101__269 clknet_1_0__leaf__02741_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__inv_2
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20202_ net262 _01133_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09944_ rbzero.tex_r0\[27\] rbzero.tex_r0\[26\] _03017_ vssd1 vssd1 vccd1 vccd1 _03025_
+ sky130_fd_sc_hd__mux2_1
X_20133_ clknet_leaf_89_i_clk _01064_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_48_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20064_ clknet_leaf_0_i_clk _00995_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09875_ rbzero.tex_r0\[60\] rbzero.tex_r0\[59\] _02984_ vssd1 vssd1 vccd1 vccd1 _02989_
+ sky130_fd_sc_hd__mux2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_1_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10650_ rbzero.map_overlay.i_mapdy\[1\] vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__inv_2
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18980__160 clknet_1_1__leaf__02729_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__inv_2
XFILLER_10_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10581_ rbzero.debug_overlay.playerX\[0\] _03373_ _03374_ rbzero.debug_overlay.playerY\[1\]
+ _03376_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__a221o_1
XFILLER_166_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12320_ _05065_ _05069_ _05071_ _05076_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__a211oi_4
XFILLER_182_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12251_ _04924_ _05008_ _05010_ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__a21o_1
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11202_ rbzero.tex_r1\[23\] _03733_ _03986_ _03666_ vssd1 vssd1 vccd1 vccd1 _03987_
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12182_ _04931_ _04943_ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__and2_1
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11133_ rbzero.tex_r1\[55\] _03618_ _03916_ _03917_ vssd1 vssd1 vccd1 vccd1 _03918_
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16990_ _09496_ _09565_ _09594_ vssd1 vssd1 vccd1 vccd1 _09596_ sky130_fd_sc_hd__and3_1
XFILLER_1_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11064_ _03834_ rbzero.map_overlay.i_mapdy\[1\] vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__xnor2_1
X_15941_ _08512_ _08558_ _08559_ _08522_ vssd1 vssd1 vccd1 vccd1 _08560_ sky130_fd_sc_hd__a31o_1
XFILLER_153_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10015_ _03062_ vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__clkbuf_1
X_18660_ _03338_ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__clkbuf_4
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15872_ rbzero.wall_tracer.mapX\[9\] _07826_ vssd1 vssd1 vccd1 vccd1 _08499_ sky130_fd_sc_hd__xnor2_1
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17611_ rbzero.debug_overlay.playerY\[0\] _03352_ _09620_ vssd1 vssd1 vccd1 vccd1
+ _01894_ sky130_fd_sc_hd__mux2_1
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14823_ _07503_ _07509_ vssd1 vssd1 vccd1 vccd1 _07511_ sky130_fd_sc_hd__and2b_1
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18591_ rbzero.pov.spi_buffer\[63\] rbzero.pov.spi_buffer\[64\] _02510_ vssd1 vssd1
+ vccd1 vccd1 _02515_ sky130_fd_sc_hd__mux2_1
XFILLER_76_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17542_ rbzero.wall_tracer.rayAddendY\[4\] rbzero.wall_tracer.rayAddendY\[3\] _01786_
+ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__o21ai_1
X_11966_ net30 net29 net31 vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__a21oi_1
XFILLER_17_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14754_ _07415_ _07441_ vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__nand2_1
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10917_ _03677_ _03695_ _03698_ _03701_ _03702_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__o221a_1
X_13705_ _06458_ _06461_ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__nand2_1
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17473_ _01764_ _01765_ _01766_ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__and3_1
X_14685_ _07361_ _07359_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__and2b_1
X_11897_ net21 vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__buf_2
XFILLER_44_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16424_ _08018_ vssd1 vssd1 vccd1 vccd1 _09035_ sky130_fd_sc_hd__clkbuf_4
X_13636_ _06349_ _06390_ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__nor2_1
XFILLER_60_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10848_ _03567_ _03603_ _03604_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__nor3_4
XFILLER_20_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19143_ clknet_1_1__leaf__02743_ vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__buf_1
XFILLER_160_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13567_ _06308_ _06323_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__xor2_1
X_16355_ rbzero.wall_tracer.trackDistX\[2\] _08553_ _08959_ _08966_ vssd1 vssd1 vccd1
+ vccd1 _00551_ sky130_fd_sc_hd__o22a_1
X_10779_ _03563_ _03564_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__or2_1
XFILLER_173_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15306_ _06997_ vssd1 vssd1 vccd1 vccd1 _07992_ sky130_fd_sc_hd__clkbuf_4
X_12518_ _05242_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__inv_2
X_16286_ _08895_ _08897_ vssd1 vssd1 vccd1 vccd1 _08898_ sky130_fd_sc_hd__xnor2_1
XFILLER_173_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13498_ _06244_ _06249_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__xor2_1
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18025_ _02214_ vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15237_ _07796_ _07923_ vssd1 vssd1 vccd1 vccd1 _07924_ sky130_fd_sc_hd__xnor2_2
X_12449_ _05153_ _05077_ _05081_ _05188_ _05205_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__o2111a_1
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15168_ _07708_ _07853_ _07854_ vssd1 vssd1 vccd1 vccd1 _07855_ sky130_fd_sc_hd__o21ai_1
XFILLER_99_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14119_ rbzero.wall_tracer.stepDistX\[-3\] _06712_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _06824_ sky130_fd_sc_hd__mux2_1
X_19976_ net205 _00907_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[56\] sky130_fd_sc_hd__dfxtp_1
X_15099_ _07786_ vssd1 vssd1 vccd1 vccd1 _07787_ sky130_fd_sc_hd__buf_2
XFILLER_80_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18858_ rbzero.pov.ready_buffer\[10\] _02635_ _02691_ _02285_ vssd1 vssd1 vccd1 vccd1
+ _01069_ sky130_fd_sc_hd__o211a_1
XFILLER_95_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17809_ _02068_ _02069_ _02072_ _02073_ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__o211ai_2
X_18789_ rbzero.pov.ready_buffer\[22\] _02644_ _02654_ _02651_ vssd1 vssd1 vccd1 vccd1
+ _01037_ sky130_fd_sc_hd__a211o_1
X_19181__341 clknet_1_1__leaf__02749_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__inv_2
XFILLER_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18904__91 clknet_1_1__leaf__02441_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__inv_2
XFILLER_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20116_ clknet_leaf_90_i_clk _01047_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[10\]
+ sky130_fd_sc_hd__dfxtp_2
X_09927_ rbzero.tex_r0\[35\] rbzero.tex_r0\[34\] _03006_ vssd1 vssd1 vccd1 vccd1 _03016_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09858_ _02978_ vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__clkbuf_1
X_20047_ clknet_leaf_81_i_clk _00978_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09789_ rbzero.tex_r1\[34\] rbzero.tex_r1\[35\] _02932_ vssd1 vssd1 vccd1 vccd1 _02942_
+ sky130_fd_sc_hd__mux2_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ net45 _04568_ _04577_ _04596_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__a31o_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ net49 _04512_ _04519_ net39 vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__a22o_1
XFILLER_42_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10702_ _03490_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__buf_4
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _04840_ rbzero.wall_tracer.stepDistX\[3\] vssd1 vssd1 vccd1 vccd1 _07158_
+ sky130_fd_sc_hd__nor2_1
X_11682_ rbzero.tex_b1\[3\] _03696_ _03697_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__and3_1
XFILLER_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13421_ _06166_ _06175_ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__nand2_1
X_10633_ _03422_ _03428_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__and2_1
X_16140_ _08742_ _08751_ vssd1 vssd1 vccd1 vccd1 _08753_ sky130_fd_sc_hd__or2_1
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13352_ _06107_ _06108_ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__nand2_1
X_10564_ rbzero.debug_overlay.playerY\[5\] vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__inv_2
XFILLER_128_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12303_ _05028_ _05029_ _05057_ _05059_ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__a31o_2
XFILLER_10_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16071_ _08680_ _07673_ _08684_ vssd1 vssd1 vccd1 vccd1 _08685_ sky130_fd_sc_hd__mux2_1
X_13283_ _06027_ _06025_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__and2b_1
X_10495_ _03314_ vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15022_ _07706_ _07707_ _07709_ vssd1 vssd1 vccd1 vccd1 _07710_ sky130_fd_sc_hd__o21ai_1
XFILLER_136_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12234_ _04961_ rbzero.wall_tracer.trackDistX\[3\] _04962_ rbzero.wall_tracer.trackDistX\[2\]
+ _04995_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__o221a_1
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19830_ clknet_leaf_4_i_clk _00761_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_mapdx\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12165_ _04881_ _04921_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__and2_2
XFILLER_64_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11116_ gpout0.vpos\[5\] vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__buf_4
X_19761_ clknet_leaf_85_i_clk _00692_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16973_ _09481_ vssd1 vssd1 vccd1 vccd1 _09579_ sky130_fd_sc_hd__inv_2
X_12096_ rbzero.debug_overlay.facingY\[-7\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__or2_1
XFILLER_111_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18712_ _06958_ _02535_ vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__nor2_1
X_11047_ _03517_ rbzero.debug_overlay.playerY\[0\] vssd1 vssd1 vccd1 vccd1 _03833_
+ sky130_fd_sc_hd__xor2_1
X_15924_ _08512_ _08543_ _08544_ _08522_ vssd1 vssd1 vccd1 vccd1 _08545_ sky130_fd_sc_hd__a31o_1
X_19692_ clknet_leaf_5_i_clk _00623_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.a6 sky130_fd_sc_hd__dfxtp_2
X_19130__295 clknet_1_1__leaf__02744_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__inv_2
XFILLER_162_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput9 i_gpout1_sel[0] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_6
XFILLER_92_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18643_ rbzero.pov.ready_buffer\[62\] _06929_ _02540_ vssd1 vssd1 vccd1 vccd1 _02547_
+ sky130_fd_sc_hd__mux2_1
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _03341_ vssd1 vssd1 vccd1 vccd1 _08485_ sky130_fd_sc_hd__buf_4
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14806_ _07039_ vssd1 vssd1 vccd1 vccd1 _07494_ sky130_fd_sc_hd__clkbuf_4
XFILLER_18_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18574_ rbzero.pov.spi_buffer\[55\] rbzero.pov.spi_buffer\[56\] _02499_ vssd1 vssd1
+ vccd1 vccd1 _02506_ sky130_fd_sc_hd__mux2_1
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15786_ rbzero.row_render.size\[2\] _08449_ _06686_ _08454_ vssd1 vssd1 vccd1 vccd1
+ _00494_ sky130_fd_sc_hd__a22o_1
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ _05752_ _05753_ _05754_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__a21oi_1
XFILLER_51_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17525_ _01784_ rbzero.wall_tracer.rayAddendY\[4\] vssd1 vssd1 vccd1 vccd1 _01815_
+ sky130_fd_sc_hd__xor2_1
XFILLER_18_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14737_ _07374_ _07424_ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__xnor2_2
X_11949_ net31 net32 vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__nor2_1
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17456_ _01746_ _01747_ _01749_ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__a21o_1
XFILLER_20_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14668_ _07008_ _06996_ vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__xnor2_1
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16407_ _09015_ _09017_ vssd1 vssd1 vccd1 vccd1 _09018_ sky130_fd_sc_hd__nand2_1
X_13619_ _06360_ _06361_ _06374_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__nand3_1
X_17387_ _03369_ _07826_ vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__xnor2_1
X_14599_ _07239_ _07263_ _07286_ vssd1 vssd1 vccd1 vccd1 _07287_ sky130_fd_sc_hd__a21o_1
XFILLER_146_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16338_ _08947_ _08948_ vssd1 vssd1 vccd1 vccd1 _08950_ sky130_fd_sc_hd__nand2_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16269_ _08879_ _08880_ vssd1 vssd1 vccd1 vccd1 _08881_ sky130_fd_sc_hd__nand2_1
XFILLER_134_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18008_ _02205_ vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19959_ net188 _00890_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1091 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19107__275 clknet_1_1__leaf__02741_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__inv_2
XFILLER_24_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_81_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_96_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10280_ rbzero.tex_b1\[59\] rbzero.tex_b1\[60\] _03199_ vssd1 vssd1 vccd1 vccd1 _03202_
+ sky130_fd_sc_hd__mux2_1
XFILLER_118_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19188__347 clknet_1_1__leaf__02750_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__inv_2
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13970_ _04836_ vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__buf_4
XFILLER_19_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12921_ _05675_ _05676_ _05677_ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__a21oi_1
XFILLER_47_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_34_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_15640_ _08201_ _08218_ _08216_ vssd1 vssd1 vccd1 vccd1 _08323_ sky130_fd_sc_hd__a21o_1
XFILLER_132_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _05392_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__buf_2
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _03911_ _04577_ _04570_ _04579_ net42 vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__a32o_1
XFILLER_27_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _08244_ _08254_ vssd1 vssd1 vccd1 vccd1 _08255_ sky130_fd_sc_hd__xnor2_1
X_12783_ _05537_ _05539_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__nand2_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17310_ rbzero.wall_tracer.trackDistY\[7\] rbzero.wall_tracer.stepDistY\[7\] vssd1
+ vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__nand2_1
XFILLER_14_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ net4 net3 vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__nor2_1
X_14522_ _07191_ _07203_ vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18290_ rbzero.spi_registers.got_new_floor _02323_ _02283_ _02377_ vssd1 vssd1 vccd1
+ vccd1 _00815_ sky130_fd_sc_hd__a31o_1
XFILLER_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_49_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17241_ _01572_ _01573_ _01574_ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__o21a_1
X_11665_ rbzero.tex_b1\[23\] rbzero.tex_b1\[22\] _03614_ vssd1 vssd1 vccd1 vccd1 _04446_
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14453_ _07117_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__buf_4
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13404_ _06073_ _06160_ _06097_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__a21oi_1
X_10616_ _03406_ _03399_ _03410_ _03411_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__or4_1
XFILLER_186_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17172_ rbzero.wall_tracer.trackDistX\[10\] rbzero.wall_tracer.stepDistX\[10\] vssd1
+ vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__or2_1
X_14384_ _07070_ _07071_ vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__nand2_1
X_11596_ _03656_ _04377_ _03669_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__o21a_1
XFILLER_127_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16123_ _08607_ _08610_ _08609_ vssd1 vssd1 vccd1 vccd1 _08736_ sky130_fd_sc_hd__a21boi_1
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13335_ _06001_ _06061_ _06060_ _06091_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__o31a_1
XFILLER_155_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10547_ rbzero.map_rom.f3 vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__clkbuf_4
XFILLER_182_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16054_ _08662_ _08667_ vssd1 vssd1 vccd1 vccd1 _08668_ sky130_fd_sc_hd__nand2_1
X_13266_ _05957_ _06006_ _06022_ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__o21a_1
X_10478_ _03305_ vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12217_ _04975_ rbzero.wall_tracer.trackDistX\[-9\] _04976_ rbzero.wall_tracer.trackDistX\[-10\]
+ _04978_ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__o221a_1
X_15005_ _07642_ _07691_ _07692_ vssd1 vssd1 vccd1 vccd1 _07693_ sky130_fd_sc_hd__a21o_1
XFILLER_124_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13197_ _05355_ _05593_ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__nor2_1
XFILLER_97_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19813_ clknet_leaf_2_i_clk _00744_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.mosi
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12148_ _04845_ _04846_ _04905_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__nand3_1
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19744_ clknet_leaf_76_i_clk _00675_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_16956_ _09476_ _09499_ _09474_ vssd1 vssd1 vccd1 vccd1 _09562_ sky130_fd_sc_hd__a21oi_1
X_12079_ net72 rbzero.wall_tracer.state\[5\] _04834_ vssd1 vssd1 vccd1 vccd1 _04842_
+ sky130_fd_sc_hd__and3_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15907_ _08527_ _08528_ _08526_ vssd1 vssd1 vccd1 vccd1 _08530_ sky130_fd_sc_hd__o21ai_1
X_19675_ clknet_leaf_81_i_clk _00606_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
X_16887_ _09484_ _09492_ vssd1 vssd1 vccd1 vccd1 _09494_ sky130_fd_sc_hd__or2_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18626_ net39 _02532_ _02262_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__o21ai_4
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15838_ rbzero.wall_tracer.mapX\[5\] _07825_ vssd1 vssd1 vccd1 vccd1 _08468_ sky130_fd_sc_hd__xor2_1
X_18557_ rbzero.pov.spi_buffer\[47\] rbzero.pov.spi_buffer\[48\] _02488_ vssd1 vssd1
+ vccd1 vccd1 _02497_ sky130_fd_sc_hd__mux2_1
X_15769_ _02901_ _03838_ _03459_ _04034_ vssd1 vssd1 vccd1 vccd1 _08443_ sky130_fd_sc_hd__and4_1
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17508_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__and2_1
XFILLER_127_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18488_ rbzero.pov.spi_buffer\[14\] rbzero.pov.spi_buffer\[15\] _02455_ vssd1 vssd1
+ vccd1 vccd1 _02461_ sky130_fd_sc_hd__mux2_1
XFILLER_36_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17439_ _04109_ rbzero.wall_tracer.rayAddendY\[-2\] vssd1 vssd1 vccd1 vccd1 _01735_
+ sky130_fd_sc_hd__nor2_1
XANTENNA_14 _06977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 rbzero.wall_tracer.visualWallDist\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_36 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20450_ net130 _01381_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[41\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_58 _06916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_69 net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19109_ clknet_1_0__leaf__02732_ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__buf_1
XFILLER_119_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20381_ net441 _01312_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11450_ _03912_ _04233_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__and2_1
XFILLER_149_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10401_ rbzero.tex_b1\[1\] rbzero.tex_b1\[2\] _02909_ vssd1 vssd1 vccd1 vccd1 _03265_
+ sky130_fd_sc_hd__mux2_1
X_11381_ rbzero.tex_g0\[31\] _04155_ _04156_ _03659_ vssd1 vssd1 vccd1 vccd1 _04165_
+ sky130_fd_sc_hd__a31o_1
XFILLER_109_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13120_ _05623_ _05876_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__or2_1
XFILLER_109_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10332_ rbzero.tex_b1\[34\] rbzero.tex_b1\[35\] _03221_ vssd1 vssd1 vccd1 vccd1 _03229_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13051_ _05558_ _05806_ _05807_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__o21ai_1
X_10263_ rbzero.tex_g0\[4\] rbzero.tex_g0\[3\] _03188_ vssd1 vssd1 vccd1 vccd1 _03193_
+ sky130_fd_sc_hd__mux2_1
XFILLER_106_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12002_ _04750_ _03913_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__nor2_1
XFILLER_133_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10194_ rbzero.tex_g0\[37\] rbzero.tex_g0\[36\] _03155_ vssd1 vssd1 vccd1 vccd1 _03157_
+ sky130_fd_sc_hd__mux2_1
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16810_ rbzero.wall_tracer.trackDistX\[6\] rbzero.wall_tracer.stepDistX\[6\] vssd1
+ vssd1 vccd1 vccd1 _09418_ sky130_fd_sc_hd__and2_1
X_17790_ _02054_ _02055_ _02042_ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__a21o_1
XFILLER_8_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16741_ _09334_ _09347_ vssd1 vssd1 vccd1 vccd1 _09349_ sky130_fd_sc_hd__or2_1
X_13953_ _05376_ _06701_ _06702_ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__o21ai_1
XFILLER_115_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12904_ _05526_ _05471_ _05518_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__or3_1
XFILLER_4_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19460_ clknet_leaf_54_i_clk _00406_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
X_16672_ _09167_ _08804_ vssd1 vssd1 vccd1 vccd1 _09281_ sky130_fd_sc_hd__or2b_1
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13884_ _06638_ _06639_ vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__nand2_1
XFILLER_62_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15623_ _08305_ _08306_ vssd1 vssd1 vccd1 vccd1 _08307_ sky130_fd_sc_hd__and2b_1
X_19391_ _02865_ _02866_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__nor2_1
X_12835_ _05467_ _05483_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__and2_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _02406_ vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__clkbuf_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _08236_ _08237_ vssd1 vssd1 vccd1 vccd1 _08238_ sky130_fd_sc_hd__nor2_1
XFILLER_43_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12766_ _05519_ _05522_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__xnor2_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _07109_ _07148_ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__or2_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _02361_ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__inv_2
X_11717_ _04487_ net65 _04493_ _04494_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__a211o_1
X_15485_ _08065_ _08169_ vssd1 vssd1 vccd1 vccd1 _08170_ sky130_fd_sc_hd__xnor2_2
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12697_ _05451_ _05453_ _05390_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17224_ rbzero.wall_tracer.trackDistY\[-5\] rbzero.wall_tracer.stepDistY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__and2_1
X_11648_ _03823_ _04428_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__or2_1
X_14436_ _07100_ _07122_ _07123_ _07121_ vssd1 vssd1 vccd1 vccd1 _07124_ sky130_fd_sc_hd__o31ai_1
XFILLER_30_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput12 i_gpout1_sel[3] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_6
XFILLER_168_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput23 i_gpout3_sel[2] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_4
Xinput34 i_gpout5_sel[1] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_6
X_17155_ _09021_ _08803_ vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__or2_1
Xinput45 i_reset_lock_a vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__buf_4
X_11579_ rbzero.tex_b0\[26\] _03617_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__and2_1
X_14367_ _06871_ _07052_ vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__nor2_1
XFILLER_6_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16106_ _08707_ _08708_ vssd1 vssd1 vccd1 vccd1 _08719_ sky130_fd_sc_hd__or2_1
XFILLER_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13318_ _06074_ _06068_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__xor2_1
X_17086_ _09657_ _09690_ vssd1 vssd1 vccd1 vccd1 _09691_ sky130_fd_sc_hd__xor2_1
Xclkbuf_1_1__f__02744_ clknet_0__02744_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02744_
+ sky130_fd_sc_hd__clkbuf_16
X_14298_ rbzero.wall_tracer.visualWallDist\[-3\] _06985_ _06906_ vssd1 vssd1 vccd1
+ vccd1 _06986_ sky130_fd_sc_hd__a21oi_1
XFILLER_157_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16037_ _08649_ _08650_ vssd1 vssd1 vccd1 vccd1 _08651_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13249_ _05959_ _05970_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__nor2_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17988_ rbzero.pov.spi_buffer\[47\] rbzero.pov.ready_buffer\[47\] _02186_ vssd1 vssd1
+ vccd1 vccd1 _02195_ sky130_fd_sc_hd__mux2_1
XFILLER_42_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19727_ clknet_leaf_94_i_clk _00658_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_16939_ _09543_ _09544_ vssd1 vssd1 vccd1 vccd1 _09545_ sky130_fd_sc_hd__xnor2_2
XFILLER_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19658_ clknet_leaf_16_i_clk _00589_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18609_ rbzero.pov.spi_buffer\[72\] rbzero.pov.spi_buffer\[73\] _02443_ vssd1 vssd1
+ vccd1 vccd1 _02524_ sky130_fd_sc_hd__mux2_1
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19589_ clknet_leaf_39_i_clk _00520_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20502_ clknet_leaf_42_i_clk _01433_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20433_ net493 _01364_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19219__376 clknet_1_1__leaf__02752_ vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__inv_2
XFILLER_106_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20364_ net424 _01295_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20295_ net355 _01226_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10950_ rbzero.tex_r0\[33\] rbzero.tex_r0\[32\] _03663_ vssd1 vssd1 vccd1 vccd1 _03736_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10881_ rbzero.tex_r0\[13\] rbzero.tex_r0\[12\] _03663_ vssd1 vssd1 vccd1 vccd1 _03667_
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ _05242_ _05240_ _05313_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__mux2_1
XFILLER_189_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12551_ _05304_ _05307_ _05269_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__a21o_1
XFILLER_196_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11502_ rbzero.tex_g1\[57\] rbzero.tex_g1\[56\] _03664_ vssd1 vssd1 vccd1 vccd1 _04285_
+ sky130_fd_sc_hd__mux2_1
XFILLER_145_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15270_ _07953_ _07955_ vssd1 vssd1 vccd1 vccd1 _07956_ sky130_fd_sc_hd__nor2_1
X_12482_ _05116_ _05199_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__nand2_1
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11433_ _04215_ _04216_ _03739_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__mux2_1
X_14221_ rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__xor2_1
XFILLER_172_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14152_ _06841_ rbzero.mapdxw\[0\] _06842_ vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__mux2_1
X_11364_ _03522_ _04031_ _04148_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__o21a_1
XFILLER_152_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10315_ rbzero.tex_b1\[42\] rbzero.tex_b1\[43\] _03210_ vssd1 vssd1 vccd1 vccd1 _03220_
+ sky130_fd_sc_hd__mux2_1
X_13103_ _05614_ _05626_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__or2b_1
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14083_ rbzero.wall_tracer.visualWallDist\[2\] _06796_ _06785_ rbzero.wall_tracer.trackDistY\[2\]
+ _06797_ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__o221a_1
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11295_ _04049_ _04076_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__or2b_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ _05789_ _05790_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__and2_1
X_17911_ rbzero.pov.spi_buffer\[10\] rbzero.pov.ready_buffer\[10\] _02153_ vssd1 vssd1
+ vccd1 vccd1 _02155_ sky130_fd_sc_hd__mux2_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10246_ rbzero.tex_g0\[12\] rbzero.tex_g0\[11\] _03177_ vssd1 vssd1 vccd1 vccd1 _03184_
+ sky130_fd_sc_hd__mux2_1
XFILLER_140_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18891_ _03520_ _02712_ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__or2_1
XFILLER_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17842_ rbzero.spi_registers.ss_buffer\[1\] _02981_ vssd1 vssd1 vccd1 vccd1 _02103_
+ sky130_fd_sc_hd__nor2_4
XFILLER_65_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10177_ rbzero.tex_g0\[45\] rbzero.tex_g0\[44\] _03144_ vssd1 vssd1 vccd1 vccd1 _03148_
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17773_ _02037_ _02038_ _02039_ vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__a21oi_1
X_14985_ rbzero.wall_tracer.visualWallDist\[-9\] _06855_ _07144_ rbzero.debug_overlay.playerY\[-9\]
+ _07146_ vssd1 vssd1 vccd1 vccd1 _07673_ sky130_fd_sc_hd__a221o_4
XFILLER_94_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19512_ clknet_leaf_61_i_clk _00458_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16724_ _09330_ _09331_ vssd1 vssd1 vccd1 vccd1 _09332_ sky130_fd_sc_hd__nor2_1
X_13936_ _06687_ vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19443_ gpout3.clk_div\[0\] net61 vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__nor2_1
X_16655_ _09161_ _09247_ _09263_ vssd1 vssd1 vccd1 vccd1 _09264_ sky130_fd_sc_hd__a21o_1
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13867_ _06588_ _06623_ vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__nor2_1
XFILLER_90_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15606_ _08162_ _08164_ vssd1 vssd1 vccd1 vccd1 _08290_ sky130_fd_sc_hd__nor2_1
XFILLER_37_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19374_ _02851_ _02852_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__xnor2_1
X_12818_ _05560_ _05537_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__nand2_1
X_16586_ _09194_ _09092_ vssd1 vssd1 vccd1 vccd1 _09196_ sky130_fd_sc_hd__or2b_1
X_13798_ _06511_ _06543_ _06553_ _06554_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__a22o_1
XFILLER_37_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18325_ rbzero.spi_registers.new_other\[9\] rbzero.spi_registers.spi_buffer\[9\]
+ _02388_ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__mux2_1
XFILLER_163_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15537_ _08188_ _08220_ vssd1 vssd1 vccd1 vccd1 _08221_ sky130_fd_sc_hd__xnor2_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12749_ _05505_ _05474_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__nor2_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18256_ _02117_ _02119_ _02121_ _02357_ vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__and4bb_1
X_15468_ _08137_ _08152_ vssd1 vssd1 vccd1 vccd1 _08153_ sky130_fd_sc_hd__xor2_1
XFILLER_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17207_ rbzero.wall_tracer.trackDistY\[-8\] _01523_ _01546_ _08532_ vssd1 vssd1 vccd1
+ vccd1 _00563_ sky130_fd_sc_hd__o22a_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14419_ _04830_ _07104_ _07106_ _03490_ vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__a211o_2
XFILLER_191_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18187_ rbzero.spi_registers.new_leak\[0\] _02310_ _02312_ _02301_ vssd1 vssd1 vccd1
+ vccd1 _00777_ sky130_fd_sc_hd__o211a_1
X_15399_ _08076_ _07976_ _08083_ vssd1 vssd1 vccd1 vccd1 _08084_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17138_ _09541_ _09637_ _09638_ _09640_ vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__a22o_1
XFILLER_116_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09960_ _03033_ vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__clkbuf_1
X_17069_ _08889_ _09256_ _09543_ _09542_ vssd1 vssd1 vccd1 vccd1 _09674_ sky130_fd_sc_hd__o31ai_1
Xclkbuf_1_1__f__02727_ clknet_0__02727_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02727_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20080_ clknet_leaf_84_i_clk _01011_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-9\]
+ sky130_fd_sc_hd__dfxtp_4
X_09891_ _02997_ vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__clkbuf_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20416_ net476 _01347_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20347_ net407 _01278_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18935__119 clknet_1_1__leaf__02725_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__inv_2
XFILLER_122_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10100_ _03107_ vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11080_ rbzero.map_overlay.i_mapdx\[1\] _03463_ _03865_ rbzero.map_overlay.i_mapdx\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__o22a_1
X_20278_ net338 _01209_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10031_ _03070_ vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_102_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14770_ _07456_ _07457_ vssd1 vssd1 vccd1 vccd1 _07458_ sky130_fd_sc_hd__nand2_1
X_11982_ net28 _04755_ _04739_ net32 vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__o211ai_1
XFILLER_44_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13721_ _06450_ _06463_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__xor2_1
XFILLER_17_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10933_ _03718_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__inv_4
XFILLER_71_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__02747_ clknet_0__02747_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02747_
+ sky130_fd_sc_hd__clkbuf_16
X_16440_ _07877_ _09046_ _09049_ vssd1 vssd1 vccd1 vccd1 _09051_ sky130_fd_sc_hd__o21ai_1
XFILLER_32_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10864_ rbzero.tex_r0\[7\] rbzero.tex_r0\[6\] _03649_ vssd1 vssd1 vccd1 vccd1 _03650_
+ sky130_fd_sc_hd__mux2_1
X_13652_ _05805_ _05987_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__nor2_1
XFILLER_182_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12603_ _05192_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__clkinv_2
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _08979_ _08980_ vssd1 vssd1 vccd1 vccd1 _08982_ sky130_fd_sc_hd__and2_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ rbzero.texV\[8\] _03580_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__xor2_1
XFILLER_24_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13583_ _06103_ _05995_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__nor2_1
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18110_ rbzero.spi_registers.got_new_other _02262_ vssd1 vssd1 vccd1 vccd1 _02263_
+ sky130_fd_sc_hd__nand2_2
XFILLER_200_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15322_ _07617_ _07646_ _07748_ _07756_ vssd1 vssd1 vccd1 vccd1 _08008_ sky130_fd_sc_hd__or4_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _05197_ _05189_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__or2b_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18041_ _02222_ vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__clkbuf_1
X_15253_ rbzero.wall_tracer.texu\[1\] _06853_ _07938_ _07939_ _03498_ vssd1 vssd1
+ vccd1 vccd1 _00476_ sky130_fd_sc_hd__o221a_1
XFILLER_126_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12465_ _05178_ _05180_ _05181_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__nand3b_1
XFILLER_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_90 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_90/HI o_rgb[21] sky130_fd_sc_hd__conb_1
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14204_ rbzero.debug_overlay.playerX\[-7\] _06887_ _04838_ vssd1 vssd1 vccd1 vccd1
+ _06892_ sky130_fd_sc_hd__a21oi_1
X_11416_ rbzero.tex_g0\[59\] rbzero.tex_g0\[58\] _04189_ vssd1 vssd1 vccd1 vccd1 _04200_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15184_ _07738_ _07852_ _07870_ vssd1 vssd1 vccd1 vccd1 _07871_ sky130_fd_sc_hd__a21o_1
XFILLER_126_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12396_ _05152_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__clkbuf_4
XFILLER_126_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11347_ rbzero.debug_overlay.playerX\[4\] _04064_ _04079_ rbzero.debug_overlay.playerX\[0\]
+ _04131_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__a221o_1
X_14135_ _06832_ vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19992_ clknet_leaf_95_i_clk _00923_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18943_ clknet_1_1__leaf__02440_ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__buf_1
X_11278_ _04060_ _04062_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__or2b_1
X_14066_ rbzero.wall_tracer.trackDistY\[-6\] _06786_ _06795_ vssd1 vssd1 vccd1 vccd1
+ _00433_ sky130_fd_sc_hd__o21a_1
X_10229_ rbzero.tex_g0\[20\] rbzero.tex_g0\[19\] _03166_ vssd1 vssd1 vccd1 vccd1 _03175_
+ sky130_fd_sc_hd__mux2_1
X_13017_ _05770_ _05773_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__xnor2_1
X_18874_ _02286_ _02703_ _04834_ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__and3b_1
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17825_ _02001_ rbzero.wall_tracer.rayAddendX\[9\] vssd1 vssd1 vccd1 vccd1 _02088_
+ sky130_fd_sc_hd__or2_1
Xhold1 rbzero.tex_r1\[40\] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_181_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17756_ _02023_ _02024_ rbzero.wall_tracer.rayAddendX\[3\] _08447_ vssd1 vssd1 vccd1
+ vccd1 _02025_ sky130_fd_sc_hd__a2bb2o_1
X_14968_ _07006_ _07174_ _07655_ vssd1 vssd1 vccd1 vccd1 _07656_ sky130_fd_sc_hd__and3b_1
XFILLER_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16707_ _09213_ _09243_ vssd1 vssd1 vccd1 vccd1 _09315_ sky130_fd_sc_hd__nand2_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13919_ _05347_ _06604_ _06671_ _05333_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__a211o_1
X_17687_ rbzero.wall_tracer.rayAddendX\[-2\] _00013_ _01957_ _01960_ vssd1 vssd1 vccd1
+ vccd1 _00629_ sky130_fd_sc_hd__o22a_1
XFILLER_63_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14899_ _07586_ vssd1 vssd1 vccd1 vccd1 _07587_ sky130_fd_sc_hd__inv_2
XFILLER_63_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19426_ rbzero.wall_tracer.rayAddendX\[-8\] _02868_ _08454_ _02882_ vssd1 vssd1 vccd1
+ vccd1 _01446_ sky130_fd_sc_hd__a22o_1
X_16638_ _09154_ _09163_ vssd1 vssd1 vccd1 vccd1 _09247_ sky130_fd_sc_hd__nand2_1
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19357_ _08439_ _02837_ _02838_ _02319_ rbzero.texV\[4\] vssd1 vssd1 vccd1 vccd1
+ _01421_ sky130_fd_sc_hd__a32o_1
X_16569_ _09175_ _09177_ vssd1 vssd1 vccd1 vccd1 _09179_ sky130_fd_sc_hd__and2_1
XFILLER_200_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18308_ _02387_ vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__clkbuf_4
X_19288_ _02777_ _02778_ _02779_ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__or3_1
XFILLER_148_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18239_ _02347_ vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20201_ net261 _01132_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20132_ clknet_leaf_89_i_clk _01063_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
X_09943_ _03024_ vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20063_ clknet_leaf_0_i_clk _00994_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_09874_ _02988_ vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__clkbuf_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10580_ rbzero.debug_overlay.playerY\[0\] _03352_ _03375_ rbzero.debug_overlay.playerY\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__a22o_1
XFILLER_194_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12250_ _04924_ _05008_ _05010_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__nand3_1
XFILLER_154_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11201_ rbzero.tex_r1\[22\] _03767_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__or2_1
XFILLER_135_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ _04932_ _04942_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__and2_1
XFILLER_162_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11132_ _03693_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__clkbuf_8
XFILLER_162_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11063_ gpout0.vpos\[5\] vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__inv_2
X_15940_ _08555_ _08556_ _08557_ vssd1 vssd1 vccd1 vccd1 _08559_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10014_ rbzero.tex_g1\[57\] rbzero.tex_g1\[58\] _03061_ vssd1 vssd1 vccd1 vccd1 _03062_
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15871_ rbzero.wall_tracer.mapX\[8\] _07826_ _08493_ _08496_ vssd1 vssd1 vccd1 vccd1
+ _08498_ sky130_fd_sc_hd__a22o_1
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17610_ _01893_ vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__clkbuf_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14822_ _07503_ _07509_ vssd1 vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__xnor2_1
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18590_ _02514_ vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17541_ _01801_ _01815_ vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__or2b_1
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _07411_ _07414_ vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__or2_1
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ net28 net29 net31 _04738_ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__a31o_1
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13704_ _06443_ _06459_ _06460_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__nand3_1
XFILLER_45_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10916_ _03606_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__buf_4
X_17472_ rbzero.debug_overlay.vplaneY\[-5\] _01743_ vssd1 vssd1 vccd1 vccd1 _01766_
+ sky130_fd_sc_hd__or2_1
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14684_ _07076_ _07371_ vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__xnor2_4
X_11896_ _03474_ _04668_ _04669_ _03464_ _04670_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__a221o_1
X_16423_ _08247_ _08245_ _08018_ _08391_ vssd1 vssd1 vccd1 vccd1 _09034_ sky130_fd_sc_hd__or4_1
X_13635_ _06346_ _06391_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__and2_1
X_10847_ rbzero.row_render.side _03631_ _03632_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__o21a_1
XFILLER_160_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16354_ _08562_ _08963_ _08965_ _08522_ vssd1 vssd1 vccd1 vccd1 _08966_ sky130_fd_sc_hd__a31o_1
X_13566_ _06309_ _06321_ _06322_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__a21oi_1
X_10778_ _03562_ _03542_ _03544_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__and3_1
X_15305_ _07969_ _07990_ vssd1 vssd1 vccd1 vccd1 _07991_ sky130_fd_sc_hd__xnor2_2
XFILLER_201_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12517_ _05273_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__buf_4
XFILLER_173_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16285_ _08108_ _08896_ vssd1 vssd1 vccd1 vccd1 _08897_ sky130_fd_sc_hd__nor2_1
XFILLER_145_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13497_ _06177_ _06179_ vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__xnor2_1
XFILLER_139_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18024_ rbzero.pov.spi_buffer\[64\] rbzero.pov.ready_buffer\[64\] _02208_ vssd1 vssd1
+ vccd1 vccd1 _02214_ sky130_fd_sc_hd__mux2_1
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15236_ _07921_ _07922_ vssd1 vssd1 vccd1 vccd1 _07923_ sky130_fd_sc_hd__nor2_1
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12448_ _05153_ _05149_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__or2_1
XFILLER_201_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15167_ _06857_ _06875_ _07235_ _06979_ vssd1 vssd1 vccd1 vccd1 _07854_ sky130_fd_sc_hd__or4_1
XFILLER_119_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12379_ _05030_ _05051_ _05054_ _05056_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__a31o_1
XFILLER_125_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14118_ _06823_ vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19975_ net204 _00906_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[55\] sky130_fd_sc_hd__dfxtp_1
X_15098_ rbzero.wall_tracer.visualWallDist\[5\] _06855_ vssd1 vssd1 vccd1 vccd1 _07786_
+ sky130_fd_sc_hd__nand2_2
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14049_ _06783_ _05004_ vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__or2_1
XFILLER_122_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18857_ _01786_ _02637_ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__or2_1
XFILLER_68_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17808_ _02054_ _02070_ _02071_ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__or3_1
X_18444__83 clknet_1_1__leaf__02439_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__inv_2
X_18788_ rbzero.debug_overlay.facingY\[-9\] _02645_ vssd1 vssd1 vccd1 vccd1 _02654_
+ sky130_fd_sc_hd__and2_1
XFILLER_94_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17739_ _01714_ _02008_ _08448_ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__a21o_1
XFILLER_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19409_ _02871_ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_165_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20115_ clknet_leaf_76_i_clk _01046_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_09926_ _03015_ vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__clkbuf_1
X_20046_ clknet_leaf_81_i_clk _00977_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_09857_ rbzero.tex_r1\[2\] rbzero.tex_r1\[3\] _02976_ vssd1 vssd1 vccd1 vccd1 _02978_
+ sky130_fd_sc_hd__mux2_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09788_ _02941_ vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__clkbuf_1
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _03910_ _04512_ _04519_ net69 vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__a22o_1
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10701_ rbzero.wall_tracer.state\[13\] vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__clkbuf_4
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ rbzero.tex_b1\[1\] rbzero.tex_b1\[0\] _03699_ vssd1 vssd1 vccd1 vccd1 _04462_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13420_ _06147_ _06153_ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__xor2_1
XFILLER_197_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10632_ rbzero.map_overlay.i_mapdx\[3\] _03413_ _03423_ _03424_ _03427_ vssd1 vssd1
+ vccd1 vccd1 _03428_ sky130_fd_sc_hd__o2111a_1
XFILLER_201_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13351_ _06087_ _06106_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__or2_1
X_10563_ rbzero.map_rom.i_row\[4\] vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__inv_2
XFILLER_155_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12302_ _05058_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__inv_2
X_16070_ _08681_ _08682_ _08683_ vssd1 vssd1 vccd1 vccd1 _08684_ sky130_fd_sc_hd__and3b_1
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10494_ rbzero.tex_b0\[22\] rbzero.tex_b0\[21\] _03313_ vssd1 vssd1 vccd1 vccd1 _03314_
+ sky130_fd_sc_hd__mux2_1
X_13282_ _05984_ _05985_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__and2_1
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15021_ _07266_ _07708_ vssd1 vssd1 vccd1 vccd1 _07709_ sky130_fd_sc_hd__nand2_1
X_12233_ _04969_ _04984_ _04991_ _04994_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__a31o_1
XFILLER_135_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12164_ _04924_ _04925_ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__and2_1
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11115_ _03834_ gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__nand2_4
X_16972_ _09447_ _09449_ _09446_ vssd1 vssd1 vccd1 vccd1 _09578_ sky130_fd_sc_hd__a21bo_1
XFILLER_150_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19760_ clknet_leaf_88_i_clk _00691_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_12095_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__or2_1
XFILLER_122_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18711_ net61 _02598_ vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__nor2_1
X_11046_ gpout0.vpos\[5\] rbzero.debug_overlay.playerY\[2\] vssd1 vssd1 vccd1 vccd1
+ _03832_ sky130_fd_sc_hd__xor2_1
X_15923_ _08540_ _08541_ _08542_ vssd1 vssd1 vccd1 vccd1 _08544_ sky130_fd_sc_hd__o21ai_1
X_19691_ clknet_leaf_5_i_clk _00622_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.b6 sky130_fd_sc_hd__dfxtp_1
XFILLER_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18642_ _02534_ _02545_ _02546_ _02356_ vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__o211a_1
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15854_ _08482_ _08467_ _08481_ vssd1 vssd1 vccd1 vccd1 _08484_ sky130_fd_sc_hd__or3_1
XFILLER_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14805_ _07488_ _07492_ vssd1 vssd1 vccd1 vccd1 _07493_ sky130_fd_sc_hd__or2b_1
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ _02505_ vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__clkbuf_1
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15785_ rbzero.row_render.size\[1\] _08449_ _06679_ _08454_ vssd1 vssd1 vccd1 vccd1
+ _00493_ sky130_fd_sc_hd__a22o_1
XFILLER_18_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12997_ _05751_ _05750_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__and2b_1
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17524_ _01786_ rbzero.wall_tracer.rayAddendY\[3\] vssd1 vssd1 vccd1 vccd1 _01814_
+ sky130_fd_sc_hd__nand2_1
XFILLER_189_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ _07409_ _07422_ _07423_ vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__a21oi_2
XFILLER_17_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11948_ _04700_ _04721_ _04722_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__o21a_2
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17455_ _01746_ _01747_ _01749_ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__nand3_1
X_14667_ _07342_ _07354_ vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__xor2_1
X_11879_ _04624_ _04652_ _04654_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__a21oi_1
X_16406_ _09016_ _08133_ _08134_ _09014_ vssd1 vssd1 vccd1 vccd1 _09017_ sky130_fd_sc_hd__o22ai_1
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13618_ _06360_ _06361_ _06374_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__a21o_1
XFILLER_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17386_ _01688_ vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__clkbuf_1
X_14598_ _07272_ _07285_ vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__xnor2_1
X_16337_ _08947_ _08948_ vssd1 vssd1 vccd1 vccd1 _08949_ sky130_fd_sc_hd__nor2_1
XFILLER_186_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13549_ _06294_ _06302_ _06303_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__and3_1
XFILLER_146_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19059__231 clknet_1_0__leaf__02737_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__inv_2
XFILLER_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16268_ _08783_ _08848_ _08878_ vssd1 vssd1 vccd1 vccd1 _08880_ sky130_fd_sc_hd__nand3_1
XFILLER_146_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18007_ rbzero.pov.spi_buffer\[56\] rbzero.pov.ready_buffer\[56\] _02197_ vssd1 vssd1
+ vccd1 vccd1 _02205_ sky130_fd_sc_hd__mux2_1
X_15219_ _07891_ _07905_ vssd1 vssd1 vccd1 vccd1 _07906_ sky130_fd_sc_hd__xnor2_2
X_16199_ _08797_ _08811_ vssd1 vssd1 vccd1 vccd1 _08812_ sky130_fd_sc_hd__xnor2_2
XFILLER_160_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_0_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19958_ net187 _00889_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19889_ clknet_leaf_24_i_clk _00820_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_110_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09909_ rbzero.tex_r0\[44\] rbzero.tex_r0\[43\] _03006_ vssd1 vssd1 vccd1 vccd1 _03007_
+ sky130_fd_sc_hd__mux2_1
XFILLER_116_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18408__50 clknet_1_0__leaf__02436_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__inv_2
XFILLER_24_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12920_ _05665_ _05674_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__nor2_1
X_20029_ clknet_leaf_85_i_clk _00960_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _05606_ _05607_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18423__64 clknet_1_0__leaf__02437_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__inv_2
XFILLER_34_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _04566_ _04577_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__and2_1
XFILLER_199_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15570_ _08251_ _08253_ vssd1 vssd1 vccd1 vccd1 _08254_ sky130_fd_sc_hd__xnor2_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12782_ _05355_ _05536_ _05538_ _05235_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14521_ _07128_ _07208_ vssd1 vssd1 vccd1 vccd1 _07209_ sky130_fd_sc_hd__xnor2_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ net4 _04509_ _04510_ net7 net8 vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__o2111a_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17240_ _01572_ _01573_ _01574_ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__nor3_1
X_14452_ _07119_ _07110_ _07137_ _07139_ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__o31a_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11664_ rbzero.tex_b1\[21\] rbzero.tex_b1\[20\] _03616_ vssd1 vssd1 vccd1 vccd1 _04445_
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13403_ _05996_ _06159_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__or2_1
X_17171_ _09711_ _09712_ _09710_ vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__a21bo_1
X_10615_ _03369_ _03358_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__nand2_1
XFILLER_128_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14383_ _07065_ _07069_ vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__xor2_1
X_11595_ rbzero.tex_b0\[5\] rbzero.tex_b0\[4\] _04376_ vssd1 vssd1 vccd1 vccd1 _04377_
+ sky130_fd_sc_hd__mux2_1
X_16122_ _08730_ _08734_ vssd1 vssd1 vccd1 vccd1 _08735_ sky130_fd_sc_hd__xnor2_1
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13334_ _06059_ _06063_ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__or2b_1
XFILLER_128_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10546_ rbzero.debug_overlay.playerX\[1\] vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__inv_2
XFILLER_10_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16053_ _08665_ _08666_ vssd1 vssd1 vccd1 vccd1 _08667_ sky130_fd_sc_hd__xnor2_1
XFILLER_109_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13265_ _06020_ _06021_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__and2_1
X_10477_ rbzero.tex_b0\[30\] rbzero.tex_b0\[29\] _03302_ vssd1 vssd1 vccd1 vccd1 _03305_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15004_ _07611_ _07641_ vssd1 vssd1 vccd1 vccd1 _07692_ sky130_fd_sc_hd__and2_1
X_12216_ _04976_ rbzero.wall_tracer.trackDistX\[-10\] _04977_ rbzero.wall_tracer.trackDistX\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__a211o_1
XFILLER_155_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13196_ _05768_ _05914_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__and2_1
XFILLER_151_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19812_ clknet_leaf_2_i_clk _00743_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.mosi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12147_ _04846_ _04905_ _04845_ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__a21o_1
XFILLER_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19743_ clknet_leaf_75_i_clk _00674_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_16955_ _09536_ _09560_ vssd1 vssd1 vccd1 vccd1 _09561_ sky130_fd_sc_hd__xor2_2
X_12078_ _04841_ _03486_ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__nor2_1
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11029_ gpout0.hpos\[4\] _03804_ _03803_ _03460_ _03814_ vssd1 vssd1 vccd1 vccd1
+ _03815_ sky130_fd_sc_hd__o221a_1
X_15906_ _08526_ _08527_ _08528_ vssd1 vssd1 vccd1 vccd1 _08529_ sky130_fd_sc_hd__or3_1
X_16886_ _09484_ _09492_ vssd1 vssd1 vccd1 vccd1 _09493_ sky130_fd_sc_hd__nand2_1
X_19674_ clknet_leaf_78_i_clk _00605_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18625_ rbzero.pov.ready _02412_ vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__and2_1
X_15837_ rbzero.map_rom.i_col\[4\] rbzero.wall_tracer.mapX\[5\] _07825_ vssd1 vssd1
+ vccd1 vccd1 _08467_ sky130_fd_sc_hd__o21a_1
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18556_ _02496_ vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__clkbuf_1
X_15768_ _04076_ _08438_ vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__nor2_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17507_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[2\] _01776_
+ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__o21bai_1
X_14719_ _07376_ _07392_ vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__or2b_1
X_18487_ _02460_ vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__clkbuf_1
X_15699_ _07581_ _07756_ _07757_ _07100_ vssd1 vssd1 vccd1 vccd1 _08382_ sky130_fd_sc_hd__o22a_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17438_ rbzero.wall_tracer.rayAddendY\[-3\] _00013_ _01731_ _01734_ vssd1 vssd1 vccd1
+ vccd1 _00606_ sky130_fd_sc_hd__o22a_1
XFILLER_178_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_15 _07052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_26 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_37 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_48 net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17369_ rbzero.spi_registers.new_mapd\[13\] rbzero.spi_registers.spi_buffer\[13\]
+ _01662_ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__mux2_1
XANTENNA_59 _06916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20380_ net440 _01311_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19113__280 clknet_1_0__leaf__02742_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__inv_2
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10400_ _03264_ vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11380_ rbzero.tex_g0\[30\] _03700_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__and2_1
XFILLER_109_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10331_ _03228_ vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10262_ _03192_ vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__clkbuf_1
X_13050_ _05494_ _05489_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__nand2_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12001_ net32 _04774_ net28 net29 vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__and4b_1
X_10193_ _03156_ vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16740_ _09334_ _09347_ vssd1 vssd1 vccd1 vccd1 _09348_ sky130_fd_sc_hd__nand2_1
XFILLER_143_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13952_ _05310_ _06666_ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__or2_1
XFILLER_19_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12903_ _05658_ _05659_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__and2b_1
XFILLER_74_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16671_ _08805_ _09167_ vssd1 vssd1 vccd1 vccd1 _09280_ sky130_fd_sc_hd__or2b_2
X_13883_ _05349_ _06623_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__or2_1
XFILLER_189_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15622_ _08303_ _08304_ vssd1 vssd1 vccd1 vccd1 _08306_ sky130_fd_sc_hd__nand2_1
X_19390_ _02860_ _02863_ _02864_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__a21oi_1
X_12834_ _05491_ _05477_ _05450_ _05479_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__and4_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ rbzero.spi_registers.new_vshift\[4\] rbzero.spi_registers.spi_buffer\[4\]
+ _02401_ vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__mux2_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _08234_ _08235_ vssd1 vssd1 vccd1 vccd1 _08237_ sky130_fd_sc_hd__and2_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12765_ _05520_ _05521_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__xor2_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _07182_ _07184_ vssd1 vssd1 vccd1 vccd1 _07192_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18272_ _02367_ vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__clkbuf_1
X_11716_ net6 net7 vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__nand2_1
X_15484_ _08166_ _08168_ vssd1 vssd1 vccd1 vccd1 _08169_ sky130_fd_sc_hd__xor2_2
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _05380_ _05385_ _05452_ _05376_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__a211o_1
XFILLER_159_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17223_ rbzero.wall_tracer.trackDistY\[-5\] rbzero.wall_tracer.stepDistY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__nor2_1
XFILLER_174_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14435_ _07092_ vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__clkbuf_4
X_11647_ rbzero.tex_b1\[55\] rbzero.tex_b1\[54\] _03615_ vssd1 vssd1 vccd1 vccd1 _04428_
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput13 i_gpout1_sel[4] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_6
XFILLER_174_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17154_ _09142_ _09110_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__nor2_1
Xinput24 i_gpout3_sel[3] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_4
Xinput35 i_gpout5_sel[2] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_6
X_14366_ _07042_ _07053_ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__xor2_1
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11578_ _04358_ _04359_ _03666_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__mux2_1
Xinput46 i_reset_lock_b vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__buf_6
X_16105_ _04966_ _08489_ _08718_ vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__a21oi_1
XFILLER_171_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13317_ _05472_ _05992_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__or2_1
X_17085_ _09658_ _09689_ vssd1 vssd1 vccd1 vccd1 _09690_ sky130_fd_sc_hd__xor2_1
Xclkbuf_1_1__f__02743_ clknet_0__02743_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02743_
+ sky130_fd_sc_hd__clkbuf_16
X_10529_ rbzero.tex_b0\[5\] rbzero.tex_b0\[4\] _03324_ vssd1 vssd1 vccd1 vccd1 _03332_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14297_ _06859_ vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__clkbuf_4
XFILLER_192_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16036_ _07281_ _07138_ vssd1 vssd1 vccd1 vccd1 _08650_ sky130_fd_sc_hd__or2_1
X_13248_ _05976_ _05974_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__and2b_1
XFILLER_69_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13179_ _05873_ _05911_ _05935_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__a21o_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_80_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_112_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17987_ _02194_ vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19726_ clknet_leaf_95_i_clk _00657_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_16938_ _08889_ _09256_ vssd1 vssd1 vccd1 vccd1 _09544_ sky130_fd_sc_hd__nor2_1
XFILLER_38_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19657_ clknet_leaf_16_i_clk _00588_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16869_ _09474_ _09475_ vssd1 vssd1 vccd1 vccd1 _09476_ sky130_fd_sc_hd__nor2_1
XFILLER_93_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_95_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18608_ _02523_ vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19588_ clknet_leaf_38_i_clk _00519_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
X_18402__45 clknet_1_1__leaf__02435_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__inv_2
XFILLER_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18539_ _02487_ vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20501_ clknet_leaf_42_i_clk _01432_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20432_ net492 _01363_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20363_ net423 _01294_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_106_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20294_ net354 _01225_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_48_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10880_ _03635_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__buf_4
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12550_ _05305_ _05302_ _05306_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__or3_1
XFILLER_12_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11501_ _04281_ _04282_ _04283_ _03726_ _03671_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__o221a_1
XFILLER_19_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12481_ _05236_ _05237_ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__xnor2_4
XFILLER_200_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14220_ _06902_ _06905_ _06906_ _06907_ vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__a2bb2o_4
X_11432_ rbzero.tex_g0\[47\] rbzero.tex_g0\[46\] _04188_ vssd1 vssd1 vccd1 vccd1 _04216_
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14151_ _03389_ _03429_ vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__and2_1
X_11363_ _03522_ _04145_ _04147_ _03910_ _03911_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__a311oi_4
XFILLER_138_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13102_ _05612_ _05613_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__or2b_1
XFILLER_180_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10314_ _03219_ vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__clkbuf_1
X_14082_ rbzero.wall_tracer.trackDistY\[1\] _06786_ _06804_ vssd1 vssd1 vccd1 vccd1
+ _00440_ sky130_fd_sc_hd__o21a_1
XFILLER_113_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11294_ _04051_ _04062_ _04060_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__nor3_4
XFILLER_65_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13033_ _05746_ _05748_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__xor2_1
X_17910_ _02154_ vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__clkbuf_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10245_ _03183_ vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18890_ _03520_ _03902_ _02260_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__and3_1
XFILLER_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10176_ _03147_ vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17841_ rbzero.spi_registers.sclk_buffer\[2\] rbzero.spi_registers.sclk_buffer\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__nor2b_2
XFILLER_191_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14984_ _06865_ vssd1 vssd1 vccd1 vccd1 _07672_ sky130_fd_sc_hd__inv_2
X_17772_ _02000_ rbzero.wall_tracer.rayAddendX\[5\] vssd1 vssd1 vccd1 vccd1 _02039_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_66_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19511_ clknet_leaf_61_i_clk _00457_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16723_ _09328_ _09329_ vssd1 vssd1 vccd1 vccd1 _09331_ sky130_fd_sc_hd__and2_1
X_13935_ rbzero.wall_tracer.stepDistY\[-6\] _06686_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _06687_ sky130_fd_sc_hd__mux2_1
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16654_ _09261_ _09262_ vssd1 vssd1 vccd1 vccd1 _09263_ sky130_fd_sc_hd__or2_1
XFILLER_35_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19442_ _02892_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__clkbuf_1
X_13866_ _06567_ _06566_ _06568_ _06622_ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__o2bb2a_1
X_15605_ _08221_ _08288_ vssd1 vssd1 vccd1 vccd1 _08289_ sky130_fd_sc_hd__xnor2_1
X_12817_ _05571_ _05572_ _05573_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__a21bo_1
X_16585_ _09092_ _09194_ vssd1 vssd1 vccd1 vccd1 _09195_ sky130_fd_sc_hd__or2b_1
X_19373_ _02844_ _02847_ _02845_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__a21boi_1
XFILLER_37_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13797_ _06530_ _06542_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__nor2_1
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15536_ _08190_ _08219_ vssd1 vssd1 vccd1 vccd1 _08220_ sky130_fd_sc_hd__xnor2_1
X_18324_ _02396_ vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__clkbuf_1
X_12748_ _05404_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__buf_2
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18255_ rbzero.spi_registers.spi_done _02244_ vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__nor2_1
X_15467_ _08150_ _08151_ vssd1 vssd1 vccd1 vccd1 _08152_ sky130_fd_sc_hd__nand2_1
X_12679_ _05367_ _05405_ _05435_ _05274_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__o211ai_1
XFILLER_187_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17206_ _01534_ _01544_ _01545_ _01527_ vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__a31o_1
XFILLER_129_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14418_ _06849_ _04915_ _07105_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1
+ _07106_ sky130_fd_sc_hd__o211a_1
X_18186_ rbzero.floor_leak\[0\] _02311_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__or2_1
X_15398_ _08080_ _08082_ vssd1 vssd1 vccd1 vccd1 _08083_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17137_ _01479_ _01480_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14349_ _04948_ _07031_ _07036_ vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__o21ai_4
XFILLER_7_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17068_ _08896_ _09110_ _09583_ _09581_ vssd1 vssd1 vccd1 vccd1 _09673_ sky130_fd_sc_hd__o31a_1
Xclkbuf_1_1__f__02726_ clknet_0__02726_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02726_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16019_ _08605_ _08606_ _08632_ vssd1 vssd1 vccd1 vccd1 _08633_ sky130_fd_sc_hd__a21o_1
X_09890_ rbzero.tex_r0\[53\] rbzero.tex_r0\[52\] _02995_ vssd1 vssd1 vccd1 vccd1 _02997_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19709_ clknet_leaf_71_i_clk _00640_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19225__381 clknet_1_1__leaf__02753_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__inv_2
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20415_ net475 _01346_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20346_ net406 _01277_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20277_ net337 _01208_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10030_ rbzero.tex_g1\[49\] rbzero.tex_g1\[50\] _03061_ vssd1 vssd1 vccd1 vccd1 _03070_
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11981_ _04507_ _04508_ _03520_ _03515_ _04750_ net29 vssd1 vssd1 vccd1 vccd1 _04755_
+ sky130_fd_sc_hd__mux4_1
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13720_ _06475_ _06476_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__nor2_1
XFILLER_17_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10932_ _03717_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__buf_6
XFILLER_44_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__02746_ clknet_0__02746_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02746_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_140_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13651_ _06122_ _05994_ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__nor2_1
X_10863_ _03615_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__buf_6
XFILLER_182_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12602_ _05357_ _05358_ _05325_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__mux2_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _08979_ _08980_ vssd1 vssd1 vccd1 vccd1 _08981_ sky130_fd_sc_hd__nor2_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _06289_ _06338_ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__or2_1
XFILLER_158_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10794_ _03574_ _03573_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__nand2_1
XFILLER_197_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _07877_ _07766_ vssd1 vssd1 vccd1 vccd1 _08007_ sky130_fd_sc_hd__or2_1
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12533_ _05257_ _05287_ _05289_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__a21o_1
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18040_ rbzero.pov.spi_buffer\[72\] rbzero.pov.ready_buffer\[72\] _02142_ vssd1 vssd1
+ vccd1 vccd1 _02222_ sky130_fd_sc_hd__mux2_1
XFILLER_185_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15252_ _07937_ _07934_ _07935_ _04832_ vssd1 vssd1 vccd1 vccd1 _07939_ sky130_fd_sc_hd__a31o_1
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12464_ _05167_ _05168_ _05174_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__o21bai_2
XFILLER_200_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_80 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_80/HI o_rgb[9] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_91 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_91/HI zeros[0] sky130_fd_sc_hd__conb_1
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14203_ _06887_ _06890_ vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__or2_1
X_11415_ rbzero.tex_g0\[57\] rbzero.tex_g0\[56\] _03700_ vssd1 vssd1 vccd1 vccd1 _04199_
+ sky130_fd_sc_hd__mux2_1
X_15183_ _07859_ _07869_ vssd1 vssd1 vccd1 vccd1 _07870_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12395_ _03489_ _05078_ _05151_ _05080_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__o31a_1
XFILLER_181_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14134_ rbzero.wall_tracer.stepDistX\[4\] _06759_ _06825_ vssd1 vssd1 vccd1 vccd1
+ _06832_ sky130_fd_sc_hd__mux2_1
XFILLER_181_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11346_ rbzero.debug_overlay.playerX\[3\] _04059_ _04090_ rbzero.debug_overlay.playerX\[-8\]
+ _04130_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__a221o_1
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19991_ clknet_leaf_95_i_clk _00922_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_19053__226 clknet_1_0__leaf__02736_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__inv_2
XFILLER_98_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14065_ rbzero.wall_tracer.visualWallDist\[-6\] _03496_ _06791_ rbzero.wall_tracer.trackDistX\[-6\]
+ _03485_ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__o221a_1
X_11277_ _04034_ _04061_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__or2_2
XFILLER_140_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13016_ _05494_ _05488_ _05771_ _05772_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__a22o_1
X_10228_ _03174_ vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18873_ _03506_ _02702_ _04499_ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__a21o_1
XFILLER_95_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17824_ rbzero.wall_tracer.rayAddendX\[8\] _00013_ _02080_ _02087_ vssd1 vssd1 vccd1
+ vccd1 _00639_ sky130_fd_sc_hd__o22a_1
XFILLER_0_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10159_ rbzero.tex_g0\[53\] rbzero.tex_g0\[52\] _03132_ vssd1 vssd1 vccd1 vccd1 _03138_
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14967_ _07048_ _07157_ vssd1 vssd1 vccd1 vccd1 _07655_ sky130_fd_sc_hd__nor2_1
X_17755_ _02020_ _02022_ _03340_ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__o21ai_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16706_ rbzero.wall_tracer.trackDistX\[5\] _08553_ _09308_ _09314_ vssd1 vssd1 vccd1
+ vccd1 _00554_ sky130_fd_sc_hd__o22a_1
XFILLER_130_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13918_ _05347_ _06626_ vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__nor2_1
X_17686_ _01722_ _01958_ _01959_ _08460_ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__a31o_1
X_14898_ _06978_ _07148_ _07554_ _07555_ vssd1 vssd1 vccd1 vccd1 _07586_ sky130_fd_sc_hd__o22a_1
X_19425_ _01921_ _01924_ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__xor2_1
X_16637_ _09138_ _09147_ _09146_ vssd1 vssd1 vccd1 vccd1 _09246_ sky130_fd_sc_hd__a21o_1
X_13849_ _06097_ _06605_ _05447_ vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__o21a_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19356_ _02834_ _02835_ _02836_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__a21o_1
X_16568_ _09175_ _09177_ vssd1 vssd1 vccd1 vccd1 _09178_ sky130_fd_sc_hd__nor2_1
XFILLER_176_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18307_ rbzero.spi_registers.spi_done _02907_ _02111_ vssd1 vssd1 vccd1 vccd1 _02387_
+ sky130_fd_sc_hd__and3_1
XFILLER_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15519_ _07865_ _07857_ _08099_ _08098_ vssd1 vssd1 vccd1 vccd1 _08203_ sky130_fd_sc_hd__o31a_1
X_16499_ _09107_ _09108_ vssd1 vssd1 vccd1 vccd1 _09109_ sky130_fd_sc_hd__xnor2_1
X_19287_ _02777_ _02778_ _02779_ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__o21ai_1
XFILLER_175_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18238_ _03338_ _02346_ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__or2_1
XFILLER_129_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18169_ rbzero.spi_registers.new_mapd\[6\] _02290_ _02302_ _02301_ vssd1 vssd1 vccd1
+ vccd1 _00769_ sky130_fd_sc_hd__o211a_1
XFILLER_172_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20200_ net260 _01131_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20131_ clknet_leaf_89_i_clk _01062_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-6\]
+ sky130_fd_sc_hd__dfxtp_2
X_09942_ rbzero.tex_r0\[28\] rbzero.tex_r0\[27\] _03017_ vssd1 vssd1 vccd1 vccd1 _03024_
+ sky130_fd_sc_hd__mux2_1
X_20062_ clknet_leaf_1_i_clk _00993_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_09873_ rbzero.tex_r0\[61\] rbzero.tex_r0\[60\] _02984_ vssd1 vssd1 vccd1 vccd1 _02988_
+ sky130_fd_sc_hd__mux2_1
XFILLER_135_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11200_ _03978_ _03980_ _03982_ _03984_ _03648_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__o221a_1
XFILLER_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12180_ _04933_ _04940_ _04941_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__o21a_1
XFILLER_150_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11131_ rbzero.tex_r1\[54\] _03767_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__or2_1
XFILLER_122_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20329_ net389 _01260_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11062_ _03518_ _03529_ _03847_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__and3_1
XFILLER_192_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10013_ _02909_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15870_ rbzero.wall_tracer.mapX\[8\] _08489_ _08488_ _08497_ vssd1 vssd1 vccd1 vccd1
+ _00535_ sky130_fd_sc_hd__a22o_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14821_ _07504_ _07507_ _07508_ vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__a21bo_1
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17540_ _01827_ _01828_ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__nand2_1
XFILLER_57_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14752_ _07438_ _07439_ vssd1 vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__or2b_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _04737_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__inv_2
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _06452_ _06457_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__xnor2_1
XFILLER_189_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10915_ rbzero.tex_r0\[18\] _03700_ _03659_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__a21o_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17471_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__nand2_1
X_14683_ _07369_ _07370_ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__nor2_2
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11895_ net23 vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__buf_2
Xclkbuf_1_0__f__02729_ clknet_0__02729_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02729_
+ sky130_fd_sc_hd__clkbuf_16
X_16422_ _08923_ _08925_ vssd1 vssd1 vccd1 vccd1 _09033_ sky130_fd_sc_hd__or2_1
X_13634_ _06001_ _06230_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__nor2_1
X_10846_ _03539_ rbzero.row_render.wall\[1\] vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__and2_1
XFILLER_60_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16353_ _08964_ vssd1 vssd1 vccd1 vccd1 _08965_ sky130_fd_sc_hd__inv_2
XFILLER_201_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13565_ _06310_ _06320_ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__nor2_1
XFILLER_73_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10777_ _03542_ _03544_ _03562_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__a21oi_1
XFILLER_160_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15304_ _07971_ _07989_ vssd1 vssd1 vccd1 vccd1 _07990_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12516_ _05272_ _05267_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__or2b_1
XFILLER_201_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16284_ _07766_ vssd1 vssd1 vccd1 vccd1 _08896_ sky130_fd_sc_hd__buf_2
XFILLER_121_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13496_ _06235_ _06252_ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__xnor2_1
XFILLER_173_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15235_ _07919_ _07920_ vssd1 vssd1 vccd1 vccd1 _07922_ sky130_fd_sc_hd__and2_1
X_18023_ _02213_ vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__clkbuf_1
X_12447_ _05077_ _05195_ _05149_ _05081_ _05153_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__a311oi_2
XFILLER_201_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15166_ _06857_ _07235_ vssd1 vssd1 vccd1 vccd1 _07853_ sky130_fd_sc_hd__nor2_1
XFILLER_5_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18918__104 clknet_1_0__leaf__02723_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__inv_2
X_12378_ _05029_ _05134_ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__nand2_1
XFILLER_5_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14117_ rbzero.wall_tracer.stepDistX\[-4\] _06705_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _06823_ sky130_fd_sc_hd__mux2_1
X_11329_ rbzero.debug_overlay.vplaneY\[10\] _04078_ _04113_ vssd1 vssd1 vccd1 vccd1
+ _04114_ sky130_fd_sc_hd__a21oi_1
X_19974_ net203 _00905_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[54\] sky130_fd_sc_hd__dfxtp_1
X_15097_ _07269_ _07334_ _07784_ vssd1 vssd1 vccd1 vccd1 _07785_ sky130_fd_sc_hd__and3b_1
XFILLER_180_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14048_ _03495_ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__inv_2
XFILLER_140_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18856_ rbzero.pov.ready_buffer\[9\] _02635_ _02690_ _02285_ vssd1 vssd1 vccd1 vccd1
+ _01068_ sky130_fd_sc_hd__o211a_1
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17807_ _02070_ _02071_ _02054_ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__o21ai_1
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18787_ rbzero.pov.ready_buffer\[43\] _02636_ _02653_ _02643_ vssd1 vssd1 vccd1 vccd1
+ _01036_ sky130_fd_sc_hd__o211a_1
X_15999_ _08611_ _08612_ vssd1 vssd1 vccd1 vccd1 _08613_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17738_ _01992_ _02007_ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17669_ _04102_ rbzero.wall_tracer.rayAddendX\[-4\] _01935_ vssd1 vssd1 vccd1 vccd1
+ _01944_ sky130_fd_sc_hd__a21o_1
X_18964__146 clknet_1_0__leaf__02727_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__inv_2
XFILLER_63_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19408_ _02334_ _02869_ _02870_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__and3_1
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19339_ rbzero.traced_texa\[2\] rbzero.texV\[2\] vssd1 vssd1 vccd1 vccd1 _02823_
+ sky130_fd_sc_hd__nand2_1
XFILLER_148_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19036__210 clknet_1_1__leaf__02735_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__inv_2
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09925_ rbzero.tex_r0\[36\] rbzero.tex_r0\[35\] _03006_ vssd1 vssd1 vccd1 vccd1 _03015_
+ sky130_fd_sc_hd__mux2_1
X_20114_ clknet_leaf_90_i_clk _01045_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_160_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20045_ clknet_leaf_82_i_clk _00976_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_09856_ _02977_ vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__clkbuf_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09787_ rbzero.tex_r1\[35\] rbzero.tex_r1\[36\] _02932_ vssd1 vssd1 vccd1 vccd1 _02941_
+ sky130_fd_sc_hd__mux2_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450__87 clknet_1_0__leaf__02441_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__inv_2
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19082__252 clknet_1_0__leaf__02739_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__inv_2
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _03489_ _03481_ _03478_ _03486_ rbzero.wall_tracer.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _00011_ sky130_fd_sc_hd__a311o_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _04459_ _04460_ _03739_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__mux2_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10631_ _03425_ _03395_ _03364_ rbzero.map_overlay.i_mapdx\[4\] _03426_ vssd1 vssd1
+ vccd1 vccd1 _03427_ sky130_fd_sc_hd__o221a_1
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13350_ _06087_ _06106_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__nand2_1
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10562_ rbzero.map_rom.c6 vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__clkbuf_4
XFILLER_10_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12301_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[9\] vssd1
+ vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__nand2_1
XFILLER_6_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13281_ _06036_ _06037_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__and2b_1
XFILLER_182_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10493_ _03143_ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__clkbuf_4
XFILLER_33_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15020_ _06874_ _06979_ vssd1 vssd1 vccd1 vccd1 _07708_ sky130_fd_sc_hd__nor2_1
X_12232_ _04962_ rbzero.wall_tracer.trackDistX\[2\] _04990_ _04992_ _04993_ vssd1
+ vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__a221o_1
XFILLER_170_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12163_ rbzero.wall_tracer.mapY\[6\] _04923_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__or2_1
XFILLER_146_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11114_ gpout0.vpos\[4\] gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__or2_2
XFILLER_190_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16971_ _09575_ _09576_ vssd1 vssd1 vccd1 vccd1 _09577_ sky130_fd_sc_hd__xor2_1
XFILLER_151_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12094_ _04852_ _04855_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__nand2_1
XFILLER_2_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18710_ _06942_ _02597_ _02587_ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__mux2_1
XFILLER_7_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15922_ _08540_ _08541_ _08542_ vssd1 vssd1 vccd1 vccd1 _08543_ sky130_fd_sc_hd__or3_1
X_11045_ _03536_ _03766_ _03830_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__mux2_1
XFILLER_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19690_ clknet_leaf_5_i_clk _00621_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.c6 sky130_fd_sc_hd__dfxtp_1
XFILLER_65_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18641_ rbzero.debug_overlay.playerX\[-7\] _02542_ vssd1 vssd1 vccd1 vccd1 _02546_
+ sky130_fd_sc_hd__or2_1
XFILLER_65_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15853_ _08467_ _08481_ _08482_ vssd1 vssd1 vccd1 vccd1 _08483_ sky130_fd_sc_hd__o21ai_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14804_ _07489_ _07490_ _07491_ vssd1 vssd1 vccd1 vccd1 _07492_ sky130_fd_sc_hd__a21bo_1
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18572_ rbzero.pov.spi_buffer\[54\] rbzero.pov.spi_buffer\[55\] _02499_ vssd1 vssd1
+ vccd1 vccd1 _02505_ sky130_fd_sc_hd__mux2_1
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996_ _05528_ _05731_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__xnor2_1
X_15784_ rbzero.row_render.size\[0\] _08449_ _06669_ _08454_ vssd1 vssd1 vccd1 vccd1
+ _00492_ sky130_fd_sc_hd__a22o_1
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ _01745_ _01801_ _01802_ _01813_ vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__a31o_1
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14735_ _07375_ _07408_ vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__nor2_1
X_11947_ net25 net26 net67 _04686_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__or4b_1
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17454_ _01748_ _01738_ _01736_ vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__a21o_1
X_14666_ _07350_ _07352_ _07353_ vssd1 vssd1 vccd1 vccd1 _07354_ sky130_fd_sc_hd__a21oi_2
XFILLER_189_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11878_ net11 _04653_ net10 vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__a21bo_1
XFILLER_33_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16405_ _08229_ vssd1 vssd1 vccd1 vccd1 _09016_ sky130_fd_sc_hd__buf_2
X_13617_ _06363_ _06372_ _06373_ vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__a21bo_1
X_10829_ _03614_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__buf_4
X_14597_ _07283_ _07284_ vssd1 vssd1 vccd1 vccd1 _07285_ sky130_fd_sc_hd__nor2_1
X_17385_ _03353_ _01687_ _08506_ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__mux2_1
XFILLER_186_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16336_ _08727_ _08824_ _08823_ vssd1 vssd1 vccd1 vccd1 _08948_ sky130_fd_sc_hd__a21oi_1
X_13548_ _06253_ _06270_ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__xnor2_1
XFILLER_71_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16267_ _08783_ _08848_ _08878_ vssd1 vssd1 vccd1 vccd1 _08879_ sky130_fd_sc_hd__a21o_1
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13479_ _06158_ _06161_ vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__nand2_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15218_ _07903_ _07904_ vssd1 vssd1 vccd1 vccd1 _07905_ sky130_fd_sc_hd__xnor2_1
X_18006_ _02204_ vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16198_ _08808_ _08810_ vssd1 vssd1 vccd1 vccd1 _08811_ sky130_fd_sc_hd__xnor2_1
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15149_ _06873_ _07332_ _07835_ vssd1 vssd1 vccd1 vccd1 _07836_ sky130_fd_sc_hd__or3b_1
XFILLER_99_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19957_ net186 _00888_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19888_ clknet_leaf_23_i_clk _00819_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_56_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18839_ rbzero.debug_overlay.vplaneY\[-8\] _02660_ vssd1 vssd1 vccd1 vccd1 _02682_
+ sky130_fd_sc_hd__or2_1
XFILLER_95_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__02439_ _02439_ vssd1 vssd1 vccd1 vccd1 clknet_0__02439_ sky130_fd_sc_hd__clkbuf_16
XFILLER_83_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_i_clk clknet_2_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_118_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09908_ _02983_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__clkbuf_4
XFILLER_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09839_ _02968_ vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__clkbuf_1
X_20028_ clknet_leaf_85_i_clk _00959_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12850_ _05301_ _05551_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__nor2_1
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ net43 _04569_ _04577_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__and3_1
XFILLER_61_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18947__130 clknet_1_1__leaf__02726_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__inv_2
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12781_ _05526_ _05515_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__xnor2_4
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _07206_ _07207_ vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__and2b_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ net4 _04496_ net6 vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__a21o_1
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19008__186 clknet_1_0__leaf__02731_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__inv_2
X_14451_ _07119_ _07138_ _07137_ _07101_ vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__o22ai_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _04442_ _04443_ _03739_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__mux2_1
XFILLER_42_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13402_ _05990_ _06071_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__nor2_1
XFILLER_70_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17170_ _01457_ _01512_ _01513_ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__o21ai_2
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10614_ rbzero.map_rom.i_col\[4\] _03390_ _03375_ rbzero.map_rom.i_row\[4\] vssd1
+ vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__or4_1
X_14382_ _06857_ _06866_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__nor2_2
X_11594_ _03615_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__buf_4
XFILLER_31_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16121_ _08732_ _08733_ vssd1 vssd1 vccd1 vccd1 _08734_ sky130_fd_sc_hd__nor2_1
XFILLER_10_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13333_ _06058_ _06089_ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10545_ rbzero.wall_tracer.state\[1\] vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__clkinv_4
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16052_ _06997_ _08130_ vssd1 vssd1 vccd1 vccd1 _08666_ sky130_fd_sc_hd__nor2_1
XFILLER_143_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13264_ _06013_ _06019_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__or2_1
X_10476_ _03304_ vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__clkbuf_1
XFILLER_157_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15003_ _07639_ _07636_ _07689_ _07690_ _07575_ vssd1 vssd1 vccd1 vccd1 _07691_ sky130_fd_sc_hd__o2111a_2
X_12215_ rbzero.wall_tracer.trackDistY\[-11\] vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__inv_2
X_18993__172 clknet_1_0__leaf__02730_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__inv_2
X_13195_ _05861_ _05919_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__nand2_1
XFILLER_155_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19811_ clknet_leaf_3_i_clk _00742_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12146_ _04888_ _04902_ _04904_ _04907_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__or4b_1
XFILLER_150_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19742_ clknet_leaf_75_i_clk _00673_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_110_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16954_ _09537_ _09559_ vssd1 vssd1 vccd1 vccd1 _09560_ sky130_fd_sc_hd__xnor2_2
X_12077_ _04840_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__buf_4
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19089__258 clknet_1_1__leaf__02740_ vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__inv_2
XFILLER_77_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11028_ _03523_ _03806_ _03804_ gpout0.hpos\[4\] _03813_ vssd1 vssd1 vccd1 vccd1
+ _03814_ sky130_fd_sc_hd__a221o_1
X_15905_ rbzero.wall_tracer.trackDistX\[-9\] rbzero.wall_tracer.stepDistX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _08528_ sky130_fd_sc_hd__and2_1
X_19673_ clknet_leaf_82_i_clk _00604_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16885_ _09490_ _09491_ vssd1 vssd1 vccd1 vccd1 _09492_ sky130_fd_sc_hd__xor2_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18624_ _02531_ vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__clkbuf_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15836_ _08466_ vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__clkbuf_1
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18555_ rbzero.pov.spi_buffer\[46\] rbzero.pov.spi_buffer\[47\] _02488_ vssd1 vssd1
+ vccd1 vccd1 _02496_ sky130_fd_sc_hd__mux2_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12979_ _05697_ _05479_ _05538_ _05477_ vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__a22o_1
X_15767_ _04035_ _08438_ vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__nor2_1
XFILLER_92_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17506_ rbzero.wall_tracer.rayAddendY\[2\] rbzero.wall_tracer.rayAddendY\[1\] _01784_
+ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__o21ai_1
X_14718_ _07404_ _07405_ vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__and2_1
XFILLER_166_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18486_ rbzero.pov.spi_buffer\[13\] rbzero.pov.spi_buffer\[14\] _02455_ vssd1 vssd1
+ vccd1 vccd1 _02460_ sky130_fd_sc_hd__mux2_1
XFILLER_75_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15698_ _07100_ _08133_ _08380_ vssd1 vssd1 vccd1 vccd1 _08381_ sky130_fd_sc_hd__nor3_1
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17437_ _01722_ _01732_ _01733_ _08460_ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__a31o_1
XFILLER_33_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14649_ _07323_ _07330_ _07335_ vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__and3_1
XANTENNA_16 _07147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_27 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_38 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17368_ _01676_ vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_49 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16319_ _08929_ _08930_ vssd1 vssd1 vccd1 vccd1 _08931_ sky130_fd_sc_hd__nor2_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17299_ _01622_ _01623_ _01624_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__o21ai_1
XFILLER_106_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19148__311 clknet_1_1__leaf__02746_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__inv_2
XFILLER_56_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19194__353 clknet_1_0__leaf__02750_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__inv_2
XFILLER_137_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10330_ rbzero.tex_b1\[35\] rbzero.tex_b1\[36\] _03221_ vssd1 vssd1 vccd1 vccd1 _03228_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10261_ rbzero.tex_g0\[5\] rbzero.tex_g0\[4\] _03188_ vssd1 vssd1 vccd1 vccd1 _03192_
+ sky130_fd_sc_hd__mux2_1
XFILLER_178_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12000_ _04750_ net65 _04737_ _04773_ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__a211o_1
X_10192_ rbzero.tex_g0\[38\] rbzero.tex_g0\[37\] _03155_ vssd1 vssd1 vccd1 vccd1 _03156_
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19014__190 clknet_1_1__leaf__02733_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__inv_2
XFILLER_120_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13951_ _05315_ _06699_ _06700_ vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__o21ai_1
XFILLER_143_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12902_ _05652_ _05647_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16670_ _09277_ _09278_ vssd1 vssd1 vccd1 vccd1 _09279_ sky130_fd_sc_hd__and2_1
XFILLER_35_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13882_ _05324_ _06617_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__or2_1
XFILLER_100_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12833_ _05484_ _05474_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__or2_1
XFILLER_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15621_ _08303_ _08304_ vssd1 vssd1 vccd1 vccd1 _08305_ sky130_fd_sc_hd__nor2_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _02405_ vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__clkbuf_1
X_15552_ _08234_ _08235_ vssd1 vssd1 vccd1 vccd1 _08236_ sky130_fd_sc_hd__nor2_1
X_12764_ _05473_ _05471_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__or2_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14503_ _07122_ _07190_ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__xnor2_1
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11715_ _04487_ _04393_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__nor2_1
X_15483_ _07968_ _08039_ _08167_ vssd1 vssd1 vccd1 vccd1 _08168_ sky130_fd_sc_hd__a21oi_2
XFILLER_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18271_ rbzero.spi_registers.spi_buffer\[5\] rbzero.spi_registers.new_sky\[5\] _02361_
+ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__mux2_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _05380_ _05379_ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__nor2_1
XFILLER_188_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17222_ rbzero.wall_tracer.trackDistY\[-6\] _01523_ _01559_ _08546_ vssd1 vssd1 vccd1
+ vccd1 _00565_ sky130_fd_sc_hd__o22a_1
X_11646_ rbzero.tex_b1\[53\] rbzero.tex_b1\[52\] _03616_ vssd1 vssd1 vccd1 vccd1 _04427_
+ sky130_fd_sc_hd__mux2_1
X_14434_ _07110_ _07118_ _07121_ vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__a21bo_1
XFILLER_128_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 i_gpout1_sel[5] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_8
X_17153_ _09547_ _01496_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__nand2_1
X_14365_ _07049_ _07052_ vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__nor2_1
Xinput25 i_gpout3_sel[4] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_8
XFILLER_196_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput36 i_gpout5_sel[3] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_6
X_11577_ rbzero.tex_b0\[31\] rbzero.tex_b0\[30\] _03732_ vssd1 vssd1 vccd1 vccd1 _04359_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput47 i_tex_in[0] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__buf_4
XFILLER_155_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13316_ _06068_ _06072_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__nand2_1
X_16104_ _08485_ _08595_ _08596_ _08507_ _08717_ vssd1 vssd1 vccd1 vccd1 _08718_ sky130_fd_sc_hd__o311a_1
X_17084_ _09687_ _09688_ vssd1 vssd1 vccd1 vccd1 _09689_ sky130_fd_sc_hd__and2_1
XFILLER_183_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10528_ _03331_ vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__02742_ clknet_0__02742_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02742_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14296_ _03491_ _06983_ vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__nand2_1
XFILLER_171_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16035_ _08366_ _08646_ _08648_ vssd1 vssd1 vccd1 vccd1 _08649_ sky130_fd_sc_hd__a21bo_1
XFILLER_143_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13247_ _05942_ _05980_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__nand2_2
XFILLER_6_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10459_ _03295_ vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13178_ _05923_ _05934_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__xor2_1
XFILLER_97_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12129_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__nand2_1
XFILLER_97_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17986_ rbzero.pov.spi_buffer\[46\] rbzero.pov.ready_buffer\[46\] _02186_ vssd1 vssd1
+ vccd1 vccd1 _02194_ sky130_fd_sc_hd__mux2_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19725_ clknet_leaf_95_i_clk _00656_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16937_ _09540_ _09541_ _09542_ vssd1 vssd1 vccd1 vccd1 _09543_ sky130_fd_sc_hd__o21ai_2
XFILLER_42_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19656_ clknet_leaf_18_i_clk _00587_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16868_ _09472_ _09473_ vssd1 vssd1 vccd1 vccd1 _09475_ sky130_fd_sc_hd__and2_1
X_18399__42 clknet_1_1__leaf__02435_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__inv_2
XFILLER_53_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18607_ rbzero.pov.spi_buffer\[71\] rbzero.pov.spi_buffer\[72\] _02443_ vssd1 vssd1
+ vccd1 vccd1 _02523_ sky130_fd_sc_hd__mux2_1
XFILLER_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15819_ rbzero.traced_texa\[0\] _08461_ _08459_ rbzero.wall_tracer.visualWallDist\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__a22o_1
X_19587_ clknet_leaf_38_i_clk _00518_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16799_ _09095_ _09300_ _09406_ vssd1 vssd1 vccd1 vccd1 _09407_ sky130_fd_sc_hd__a21oi_1
X_18538_ rbzero.pov.spi_buffer\[38\] rbzero.pov.spi_buffer\[39\] _02477_ vssd1 vssd1
+ vccd1 vccd1 _02487_ sky130_fd_sc_hd__mux2_1
XFILLER_178_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18469_ rbzero.pov.spi_buffer\[5\] rbzero.pov.spi_buffer\[6\] _02444_ vssd1 vssd1
+ vccd1 vccd1 _02451_ sky130_fd_sc_hd__mux2_1
XFILLER_61_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20500_ clknet_leaf_42_i_clk _01431_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20431_ net491 _01362_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20362_ net422 _01293_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20293_ net353 _01224_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11500_ rbzero.tex_g1\[61\] rbzero.tex_g1\[60\] _03618_ vssd1 vssd1 vccd1 vccd1 _04283_
+ sky130_fd_sc_hd__mux2_1
XFILLER_200_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19202__360 clknet_1_0__leaf__02751_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__inv_2
XFILLER_157_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12480_ _05114_ _05119_ _05199_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__o21a_1
XFILLER_138_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ rbzero.tex_g0\[45\] rbzero.tex_g0\[44\] _04188_ vssd1 vssd1 vccd1 vccd1 _04215_
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14150_ rbzero.mapdyw\[0\] _06839_ _06840_ _03409_ vssd1 vssd1 vccd1 vccd1 _06841_
+ sky130_fd_sc_hd__a22o_1
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11362_ _03467_ _03502_ _03525_ _04146_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__or4_1
XFILLER_152_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13101_ _05630_ _05643_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__or2b_1
X_10313_ rbzero.tex_b1\[43\] rbzero.tex_b1\[44\] _03210_ vssd1 vssd1 vccd1 vccd1 _03219_
+ sky130_fd_sc_hd__mux2_1
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_1_0_i_clk clknet_1_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_152_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14081_ rbzero.wall_tracer.visualWallDist\[1\] _06796_ _06791_ rbzero.wall_tracer.trackDistX\[1\]
+ _06797_ vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__o221a_1
X_11293_ _04059_ _04069_ _04077_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__or3b_4
XFILLER_106_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13032_ _05774_ _05787_ _05788_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__a21bo_1
XFILLER_79_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10244_ rbzero.tex_g0\[13\] rbzero.tex_g0\[12\] _03177_ vssd1 vssd1 vccd1 vccd1 _03183_
+ sky130_fd_sc_hd__mux2_1
XFILLER_105_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17840_ rbzero.wall_tracer.rayAddendX\[10\] _08449_ _02101_ vssd1 vssd1 vccd1 vccd1
+ _00641_ sky130_fd_sc_hd__a21o_1
XFILLER_79_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10175_ rbzero.tex_g0\[46\] rbzero.tex_g0\[45\] _03144_ vssd1 vssd1 vccd1 vccd1 _03147_
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17771_ rbzero.wall_tracer.rayAddendX\[4\] rbzero.wall_tracer.rayAddendX\[3\] _02001_
+ vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__o21ai_1
X_14983_ _07049_ _07670_ vssd1 vssd1 vccd1 vccd1 _07671_ sky130_fd_sc_hd__nor2_1
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19510_ clknet_leaf_58_i_clk _00456_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16722_ _09328_ _09329_ vssd1 vssd1 vccd1 vccd1 _09330_ sky130_fd_sc_hd__nor2_1
XFILLER_47_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13934_ _06682_ _06685_ vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__or2_1
XFILLER_74_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19441_ _02334_ _02890_ _02891_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__and3_1
X_16653_ _09252_ _09260_ vssd1 vssd1 vccd1 vccd1 _09262_ sky130_fd_sc_hd__nor2_1
X_13865_ _06333_ _06566_ vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__nor2_1
XFILLER_170_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15604_ _08286_ _08287_ vssd1 vssd1 vccd1 vccd1 _08288_ sky130_fd_sc_hd__xor2_1
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19372_ _02849_ _02850_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__and2b_1
X_12816_ _05570_ _05555_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__or2b_1
X_16584_ _09191_ _09193_ vssd1 vssd1 vccd1 vccd1 _09194_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13796_ _06539_ _06540_ _06552_ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__a21oi_1
XFILLER_188_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18323_ rbzero.spi_registers.new_other\[8\] rbzero.spi_registers.spi_buffer\[8\]
+ _02388_ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__mux2_1
X_15535_ _08201_ _08218_ vssd1 vssd1 vccd1 vccd1 _08219_ sky130_fd_sc_hd__xor2_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12747_ _05473_ _05503_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__nor2_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18254_ rbzero.spi_registers.new_vshift\[5\] _02348_ _02355_ _02356_ vssd1 vssd1
+ vccd1 vccd1 _00800_ sky130_fd_sc_hd__o211a_1
XFILLER_179_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15466_ _08147_ _08148_ _08149_ vssd1 vssd1 vccd1 vccd1 _08151_ sky130_fd_sc_hd__o21ai_1
X_12678_ _05340_ _05341_ _05325_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__a21o_1
XFILLER_129_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17205_ _01541_ _01542_ _01543_ vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__a21o_1
X_11629_ _03612_ _04407_ _04409_ _03689_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__o211a_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14417_ _06849_ _05137_ vssd1 vssd1 vccd1 vccd1 _07105_ sky130_fd_sc_hd__nand2_1
X_18185_ rbzero.spi_registers.got_new_leak _02262_ vssd1 vssd1 vccd1 vccd1 _02311_
+ sky130_fd_sc_hd__and2_1
X_15397_ _07265_ _08081_ vssd1 vssd1 vccd1 vccd1 _08082_ sky130_fd_sc_hd__nor2_1
XFILLER_129_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17136_ _08862_ _08333_ _09663_ _09662_ _09661_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__o32a_1
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14348_ _04839_ _07035_ vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__or2_1
XFILLER_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17067_ _09670_ _09671_ vssd1 vssd1 vccd1 vccd1 _09672_ sky130_fd_sc_hd__xnor2_2
XFILLER_171_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__02725_ clknet_0__02725_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02725_
+ sky130_fd_sc_hd__clkbuf_16
X_14279_ _06940_ _06955_ _06966_ vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__or3_1
X_16018_ _08615_ _08631_ vssd1 vssd1 vccd1 vccd1 _08632_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19030__205 clknet_1_0__leaf__02734_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__inv_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ rbzero.pov.spi_buffer\[38\] rbzero.pov.ready_buffer\[38\] _02175_ vssd1 vssd1
+ vccd1 vccd1 _02185_ sky130_fd_sc_hd__mux2_1
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19708_ clknet_leaf_71_i_clk _00639_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19639_ clknet_leaf_39_i_clk _00570_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20414_ net474 _01345_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20345_ net405 _01276_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20276_ net336 _01207_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11980_ _03852_ _04750_ net29 _04753_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__a211o_1
XFILLER_99_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10931_ _03603_ _03715_ _03716_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__or3_1
XFILLER_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__02745_ clknet_0__02745_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02745_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_147_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10862_ _03627_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__buf_4
X_13650_ _05805_ _06061_ _06367_ _06369_ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__o22ai_1
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12601_ _05189_ _05197_ _05313_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__mux2_1
X_19126__291 clknet_1_0__leaf__02744_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__inv_2
XFILLER_13_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13581_ _05862_ _05992_ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__nor2_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ rbzero.texV\[7\] _03577_ _03578_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__nand3_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15320_ _08004_ _08005_ vssd1 vssd1 vccd1 vccd1 _08006_ sky130_fd_sc_hd__and2_1
XFILLER_13_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12532_ _05158_ _05175_ _05182_ _05184_ _05288_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__a41o_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12463_ _05212_ _05215_ _05217_ _05219_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__or4b_1
XFILLER_71_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15251_ _07934_ _07935_ _07937_ vssd1 vssd1 vccd1 vccd1 _07938_ sky130_fd_sc_hd__a21oi_1
XFILLER_166_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_81 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_81/HI o_rgb[10] sky130_fd_sc_hd__conb_1
X_11414_ _03607_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__buf_4
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14202_ _06888_ _06889_ vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__nand2_1
Xtop_ew_algofoogle_92 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_92/HI zeros[1] sky130_fd_sc_hd__conb_1
X_15182_ _07867_ _07868_ vssd1 vssd1 vccd1 vccd1 _07869_ sky130_fd_sc_hd__and2b_1
XFILLER_123_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12394_ rbzero.wall_tracer.visualWallDist\[10\] _03480_ vssd1 vssd1 vccd1 vccd1 _05151_
+ sky130_fd_sc_hd__nor2_1
XFILLER_125_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14133_ _06831_ vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11345_ rbzero.debug_overlay.playerX\[-9\] _04081_ _04089_ rbzero.debug_overlay.playerX\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__a22o_1
XFILLER_125_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19990_ clknet_leaf_95_i_clk _00921_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_94_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_14064_ rbzero.wall_tracer.trackDistY\[-7\] _06786_ _06794_ vssd1 vssd1 vccd1 vccd1
+ _00432_ sky130_fd_sc_hd__o21a_1
X_11276_ gpout0.hpos\[5\] _04053_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__nor2_1
XFILLER_98_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13015_ _05484_ _05489_ _05505_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__mux2_1
X_10227_ rbzero.tex_g0\[21\] rbzero.tex_g0\[20\] _03166_ vssd1 vssd1 vccd1 vccd1 _03174_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__02441_ clknet_0__02441_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02441_
+ sky130_fd_sc_hd__clkbuf_16
X_18872_ _03906_ _03531_ _02696_ _03909_ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__or4b_1
X_17823_ _01722_ _02085_ _02086_ _08460_ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__a31o_1
X_10158_ _03137_ vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17754_ _02020_ _02022_ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__and2_1
X_10089_ _03101_ vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__clkbuf_1
X_14966_ _06872_ _07148_ vssd1 vssd1 vccd1 vccd1 _07654_ sky130_fd_sc_hd__nor2_1
XFILLER_75_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16705_ _08562_ _09312_ _09313_ _08487_ vssd1 vssd1 vccd1 vccd1 _09314_ sky130_fd_sc_hd__a31o_1
X_13917_ _06670_ vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__clkbuf_1
X_17685_ rbzero.debug_overlay.vplaneX\[-6\] _01948_ vssd1 vssd1 vccd1 vccd1 _01959_
+ sky130_fd_sc_hd__or2_1
XFILLER_47_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14897_ _07552_ _07558_ vssd1 vssd1 vccd1 vccd1 _07585_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_32_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19424_ rbzero.wall_tracer.rayAddendX\[-9\] _08449_ _02881_ vssd1 vssd1 vccd1 vccd1
+ _01445_ sky130_fd_sc_hd__a21o_1
X_16636_ _09211_ _09244_ vssd1 vssd1 vccd1 vccd1 _09245_ sky130_fd_sc_hd__xnor2_1
X_13848_ _06601_ _06595_ _06597_ vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__and3_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19355_ _02834_ _02835_ _02836_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__nand3_1
X_16567_ _09030_ _09060_ _09176_ vssd1 vssd1 vccd1 vccd1 _09177_ sky130_fd_sc_hd__a21oi_1
XFILLER_188_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13779_ _06533_ _06535_ vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__xor2_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18306_ rbzero.spi_registers.got_new_leak _02323_ _02283_ _02386_ vssd1 vssd1 vccd1
+ vccd1 _00822_ sky130_fd_sc_hd__a31o_1
XFILLER_176_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15518_ _08080_ _08082_ _08079_ vssd1 vssd1 vccd1 vccd1 _08202_ sky130_fd_sc_hd__a21bo_1
XFILLER_148_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19286_ _02772_ _02775_ _02773_ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__a21boi_1
X_16498_ _07865_ _08317_ vssd1 vssd1 vccd1 vccd1 _09108_ sky130_fd_sc_hd__and2_1
XFILLER_175_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_47_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18237_ rbzero.color_floor\[5\] rbzero.spi_registers.new_floor\[5\] _02335_ vssd1
+ vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__mux2_1
X_15449_ _07757_ vssd1 vssd1 vccd1 vccd1 _08134_ sky130_fd_sc_hd__buf_2
XFILLER_30_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18168_ rbzero.map_overlay.i_mapdy\[2\] _02292_ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__or2_1
XFILLER_11_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17119_ _09636_ _01462_ _09651_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__o21ba_1
XFILLER_128_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18099_ _02254_ vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20130_ clknet_leaf_78_i_clk _01061_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-7\]
+ sky130_fd_sc_hd__dfxtp_2
X_09941_ _03023_ vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__02739_ _02739_ vssd1 vssd1 vccd1 vccd1 clknet_0__02739_ sky130_fd_sc_hd__clkbuf_16
X_20061_ clknet_leaf_1_i_clk _00992_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ss_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_09872_ _02987_ vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__clkbuf_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18941__125 clknet_1_0__leaf__02725_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__inv_2
XFILLER_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11130_ rbzero.color_sky\[1\] _03535_ _03914_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__o21ai_1
X_20328_ net388 _01259_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11061_ _03837_ _03844_ _03846_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__or3_2
X_20259_ net319 _01190_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10012_ _03060_ vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ _07451_ _07505_ vssd1 vssd1 vccd1 vccd1 _07508_ sky130_fd_sc_hd__nand2_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14751_ _07432_ _07428_ vssd1 vssd1 vccd1 vccd1 _07439_ sky130_fd_sc_hd__xnor2_1
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11963_ net30 net31 vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__nand2_1
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _06440_ _06441_ _06442_ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__a21o_1
X_10914_ _03699_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__buf_4
X_17470_ _01762_ _01763_ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__nand2_1
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14682_ _07339_ _07368_ vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__and2_1
X_11894_ net22 net21 vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_0__f__02728_ clknet_0__02728_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02728_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16421_ _07662_ _08803_ _08799_ vssd1 vssd1 vccd1 vccd1 _09032_ sky130_fd_sc_hd__or3_1
X_10845_ _03606_ _03611_ _03621_ _03630_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__a31o_1
X_13633_ _06345_ _06348_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__and2_1
XFILLER_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16352_ _08960_ _08961_ _08962_ vssd1 vssd1 vccd1 vccd1 _08964_ sky130_fd_sc_hd__and3_1
X_10776_ rbzero.texV\[5\] _03561_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__xnor2_1
X_13564_ _06310_ _06320_ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__xor2_1
XFILLER_160_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15303_ _07987_ _07988_ vssd1 vssd1 vccd1 vccd1 _07989_ sky130_fd_sc_hd__and2_1
XFILLER_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12515_ _05120_ _05243_ _05234_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__a21oi_1
X_16283_ _08892_ _08894_ vssd1 vssd1 vccd1 vccd1 _08895_ sky130_fd_sc_hd__and2_1
XFILLER_158_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13495_ _06237_ _06251_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__xor2_1
XFILLER_201_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18022_ rbzero.pov.spi_buffer\[63\] rbzero.pov.ready_buffer\[63\] _02208_ vssd1 vssd1
+ vccd1 vccd1 _02213_ sky130_fd_sc_hd__mux2_1
X_15234_ _07919_ _07920_ vssd1 vssd1 vccd1 vccd1 _07921_ sky130_fd_sc_hd__nor2_1
X_12446_ _05153_ _05077_ _05149_ _05188_ vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__o211ai_2
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15165_ _07740_ _07728_ vssd1 vssd1 vccd1 vccd1 _07852_ sky130_fd_sc_hd__or2b_1
X_12377_ rbzero.debug_overlay.facingX\[0\] rbzero.wall_tracer.rayAddendX\[8\] vssd1
+ vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__nand2_1
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11328_ rbzero.debug_overlay.vplaneY\[0\] _04079_ _04108_ _04112_ vssd1 vssd1 vccd1
+ vccd1 _04113_ sky130_fd_sc_hd__a211o_1
X_14116_ _06822_ vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__clkbuf_1
X_19973_ net202 _00904_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[53\] sky130_fd_sc_hd__dfxtp_1
X_15096_ rbzero.wall_tracer.visualWallDist\[5\] _07256_ vssd1 vssd1 vccd1 vccd1 _07784_
+ sky130_fd_sc_hd__and2_1
XFILLER_99_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11259_ _04041_ _04043_ _04035_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__or3b_1
X_14047_ _06782_ vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18855_ _01871_ _02635_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__nand2_1
XFILLER_80_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17806_ _02000_ rbzero.debug_overlay.vplaneX\[-1\] vssd1 vssd1 vccd1 vccd1 _02071_
+ sky130_fd_sc_hd__and2_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18786_ rbzero.debug_overlay.facingX\[10\] _02638_ vssd1 vssd1 vccd1 vccd1 _02653_
+ sky130_fd_sc_hd__or2_1
X_15998_ _08209_ _08325_ _08327_ _08193_ vssd1 vssd1 vccd1 vccd1 _08612_ sky130_fd_sc_hd__a22oi_2
XFILLER_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17737_ _02005_ _02006_ vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14949_ _07614_ _07635_ vssd1 vssd1 vccd1 vccd1 _07637_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19142__306 clknet_1_1__leaf__02745_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__inv_2
X_17668_ rbzero.debug_overlay.vplaneX\[-3\] rbzero.wall_tracer.rayAddendX\[-3\] vssd1
+ vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__and2_1
XFILLER_39_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19407_ gpout0.clk_div\[0\] gpout0.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__or2_1
X_16619_ _09135_ _09137_ _09134_ vssd1 vssd1 vccd1 vccd1 _09228_ sky130_fd_sc_hd__a21bo_1
X_17599_ _01858_ _01867_ _01883_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__o21ai_1
XFILLER_50_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19338_ rbzero.traced_texa\[2\] rbzero.texV\[2\] vssd1 vssd1 vccd1 vccd1 _02822_
+ sky130_fd_sc_hd__or2_1
XFILLER_176_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19269_ _02760_ _02763_ _02764_ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__nand3b_1
XFILLER_191_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20113_ clknet_leaf_90_i_clk _01044_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09924_ _03014_ vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20044_ clknet_leaf_82_i_clk _00975_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_09855_ rbzero.tex_r1\[3\] rbzero.tex_r1\[4\] _02976_ vssd1 vssd1 vccd1 vccd1 _02977_
+ sky130_fd_sc_hd__mux2_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09786_ _02940_ vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_i_clk clknet_2_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10630_ rbzero.map_overlay.i_mapdx\[1\] _03343_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__xnor2_1
XFILLER_198_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10561_ rbzero.debug_overlay.playerY\[1\] vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__inv_2
XFILLER_182_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12300_ _05030_ _05051_ _05054_ _05055_ _05056_ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__a311o_1
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13280_ _06008_ _05992_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__nor2_1
X_10492_ _03312_ vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12231_ rbzero.wall_tracer.trackDistY\[1\] rbzero.wall_tracer.trackDistX\[1\] vssd1
+ vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__and2b_1
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12162_ rbzero.wall_tracer.mapY\[6\] _04923_ vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__nand2_1
XFILLER_146_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11113_ _03534_ _03831_ _03898_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__o21a_1
X_16970_ _07993_ _08317_ vssd1 vssd1 vccd1 vccd1 _09576_ sky130_fd_sc_hd__and2_1
XFILLER_2_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12093_ _04853_ _04854_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__and2b_1
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11044_ rbzero.row_render.vinf _03822_ _03829_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__o21a_2
X_15921_ _08533_ _08535_ _08534_ vssd1 vssd1 vccd1 vccd1 _08542_ sky130_fd_sc_hd__a21boi_1
XFILLER_89_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18640_ rbzero.pov.ready_buffer\[61\] _06890_ _02540_ vssd1 vssd1 vccd1 vccd1 _02545_
+ sky130_fd_sc_hd__mux2_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15852_ rbzero.wall_tracer.mapX\[6\] _07825_ vssd1 vssd1 vccd1 vccd1 _08482_ sky130_fd_sc_hd__xor2_1
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ _06871_ _06949_ _07435_ vssd1 vssd1 vccd1 vccd1 _07491_ sky130_fd_sc_hd__or3_1
XFILLER_188_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18571_ _02504_ vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__clkbuf_1
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15783_ _08452_ vssd1 vssd1 vccd1 vccd1 _08454_ sky130_fd_sc_hd__buf_4
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12995_ _05750_ _05751_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ _01722_ _01811_ _01812_ _08448_ rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__a32o_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14734_ _07415_ _07421_ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__xnor2_1
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11946_ _04703_ _04705_ _04708_ _04720_ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__a31o_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17453_ rbzero.debug_overlay.vplaneY\[-2\] rbzero.wall_tracer.rayAddendY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__or2_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14665_ _07343_ _07349_ vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__nor2_1
XFILLER_189_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11877_ _03906_ _04499_ _03909_ _04500_ _04616_ _04612_ vssd1 vssd1 vccd1 vccd1 _04653_
+ sky130_fd_sc_hd__mux4_1
XFILLER_60_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16404_ _09014_ _08229_ _08133_ _08134_ vssd1 vssd1 vccd1 vccd1 _09015_ sky130_fd_sc_hd__or4_1
XFILLER_60_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13616_ _06364_ _06365_ _06371_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__nand3_1
X_10828_ _03556_ _03613_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__nand2_4
X_17384_ rbzero.debug_overlay.playerX\[2\] _01686_ _09620_ vssd1 vssd1 vccd1 vccd1
+ _01687_ sky130_fd_sc_hd__mux2_1
X_14596_ _07280_ _07282_ vssd1 vssd1 vccd1 vccd1 _07284_ sky130_fd_sc_hd__and2_1
XFILLER_186_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16335_ _08846_ _08946_ vssd1 vssd1 vccd1 vccd1 _08947_ sky130_fd_sc_hd__xnor2_1
XFILLER_186_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13547_ _06294_ _06302_ _06303_ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__a21oi_2
X_10759_ _03542_ _03543_ rbzero.texV\[4\] vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__a21o_1
XFILLER_173_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19054_ clknet_1_0__leaf__02732_ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__buf_1
X_16266_ _08860_ _08877_ vssd1 vssd1 vccd1 vccd1 _08878_ sky130_fd_sc_hd__xnor2_1
XFILLER_199_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13478_ _06232_ _06234_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__nand2_1
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18005_ rbzero.pov.spi_buffer\[55\] rbzero.pov.ready_buffer\[55\] _02197_ vssd1 vssd1
+ vccd1 vccd1 _02204_ sky130_fd_sc_hd__mux2_1
X_15217_ _07749_ _07759_ _07755_ vssd1 vssd1 vccd1 vccd1 _07904_ sky130_fd_sc_hd__o21a_1
XFILLER_195_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12429_ _05071_ _05076_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__nor2_1
X_16197_ _08676_ _08686_ _08809_ vssd1 vssd1 vccd1 vccd1 _08810_ sky130_fd_sc_hd__a21o_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15148_ _07049_ _07786_ vssd1 vssd1 vccd1 vccd1 _07835_ sky130_fd_sc_hd__nor2_1
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19956_ net185 _00887_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[36\] sky130_fd_sc_hd__dfxtp_1
X_15079_ _07213_ _07766_ _07180_ vssd1 vssd1 vccd1 vccd1 _07767_ sky130_fd_sc_hd__o21ba_1
XFILLER_45_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18970__151 clknet_1_1__leaf__02728_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__inv_2
XFILLER_141_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19887_ clknet_leaf_24_i_clk _00818_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18838_ rbzero.pov.ready_buffer\[0\] _02663_ _02681_ _02672_ vssd1 vssd1 vccd1 vccd1
+ _01059_ sky130_fd_sc_hd__o211a_1
XFILLER_28_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__02438_ _02438_ vssd1 vssd1 vccd1 vccd1 clknet_0__02438_ sky130_fd_sc_hd__clkbuf_16
X_18769_ _04828_ vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__buf_2
X_19066__237 clknet_1_1__leaf__02738_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__inv_2
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09907_ _03005_ vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20027_ clknet_leaf_86_i_clk _00958_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_09838_ rbzero.tex_r1\[11\] rbzero.tex_r1\[12\] _02965_ vssd1 vssd1 vccd1 vccd1 _02968_
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09769_ _02931_ vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ net18 net17 vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__nor2_2
XFILLER_55_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12780_ _05301_ _05354_ _05535_ _05536_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__or4_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _04507_ _04508_ _03520_ _03515_ _04487_ _04496_ vssd1 vssd1 vccd1 vccd1 _04509_
+ sky130_fd_sc_hd__mux4_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14450_ _07109_ vssd1 vssd1 vccd1 vccd1 _07138_ sky130_fd_sc_hd__buf_2
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ rbzero.tex_b1\[19\] rbzero.tex_b1\[18\] _03699_ vssd1 vssd1 vccd1 vccd1 _04443_
+ sky130_fd_sc_hd__mux2_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _06072_ _06157_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__nand2_1
X_10613_ _03353_ _03345_ _03394_ _03408_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__a31o_1
X_11593_ _03652_ _04374_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__or2_1
X_14381_ _07066_ _07067_ _07068_ vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__o21a_1
XFILLER_70_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16120_ _07865_ _07959_ _08070_ _07972_ vssd1 vssd1 vccd1 vccd1 _08733_ sky130_fd_sc_hd__o22a_1
XFILLER_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13332_ _06087_ _06088_ vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__xor2_1
X_10544_ _03339_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__buf_4
XFILLER_155_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16051_ _08663_ _08664_ vssd1 vssd1 vccd1 vccd1 _08665_ sky130_fd_sc_hd__nand2_1
XFILLER_183_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10475_ rbzero.tex_b0\[31\] rbzero.tex_b0\[30\] _03302_ vssd1 vssd1 vccd1 vccd1 _03304_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13263_ _06013_ _06019_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__nand2_1
XFILLER_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15002_ _07639_ _07636_ _07576_ _07608_ vssd1 vssd1 vccd1 vccd1 _07690_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19171__332 clknet_1_0__leaf__02748_ vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__inv_2
X_12214_ rbzero.wall_tracer.trackDistY\[-10\] vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__inv_2
X_13194_ _05923_ _05934_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__or2b_1
XFILLER_68_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12145_ _04905_ _04906_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__nand2_1
X_19810_ clknet_leaf_15_i_clk _00741_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16953_ _09539_ _09558_ vssd1 vssd1 vccd1 vccd1 _09559_ sky130_fd_sc_hd__xnor2_1
XFILLER_173_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19741_ clknet_leaf_75_i_clk _00672_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_12076_ _04839_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__clkbuf_4
XFILLER_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15904_ rbzero.wall_tracer.trackDistX\[-9\] rbzero.wall_tracer.stepDistX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _08527_ sky130_fd_sc_hd__nor2_1
X_11027_ gpout0.hpos\[3\] _03806_ _03808_ _03526_ _03812_ vssd1 vssd1 vccd1 vccd1
+ _03813_ sky130_fd_sc_hd__o221a_1
X_19672_ clknet_leaf_35_i_clk _00603_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16884_ _09021_ _09039_ _09364_ _09362_ vssd1 vssd1 vccd1 vccd1 _09491_ sky130_fd_sc_hd__o31a_1
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18623_ rbzero.pov.sclk_buffer\[2\] rbzero.pov.sclk_buffer\[1\] _04827_ vssd1 vssd1
+ vccd1 vccd1 _02531_ sky130_fd_sc_hd__mux2_1
XFILLER_64_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15835_ rbzero.wall_tracer.wall\[1\] rbzero.row_render.wall\[1\] _08464_ vssd1 vssd1
+ vccd1 vccd1 _08466_ sky130_fd_sc_hd__mux2_1
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18554_ _02495_ vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15766_ _04062_ _08438_ vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__nor2_1
X_12978_ _05484_ _05536_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__nor2_1
XFILLER_75_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ rbzero.wall_tracer.rayAddendY\[2\] _00013_ _01789_ _01796_ vssd1 vssd1 vccd1
+ vccd1 _00611_ sky130_fd_sc_hd__o22a_1
XFILLER_45_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14717_ _07395_ _07399_ _07403_ vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__nand3_1
X_18485_ _02459_ vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__clkbuf_1
X_11929_ _04672_ _04393_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__nor2_1
X_15697_ _07581_ _07757_ vssd1 vssd1 vccd1 vccd1 _08380_ sky130_fd_sc_hd__or2_1
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17436_ rbzero.debug_overlay.vplaneY\[-7\] _01723_ vssd1 vssd1 vccd1 vccd1 _01733_
+ sky130_fd_sc_hd__nand2_1
XFILLER_82_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14648_ _07323_ _07330_ _07335_ vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__a21oi_4
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 _07817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_28 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ rbzero.spi_registers.new_mapd\[12\] rbzero.spi_registers.spi_buffer\[12\]
+ _01662_ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__mux2_1
X_14579_ _07012_ _07265_ _07266_ vssd1 vssd1 vccd1 vccd1 _07267_ sky130_fd_sc_hd__o21bai_1
XFILLER_158_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16318_ _08927_ _08928_ vssd1 vssd1 vccd1 vccd1 _08930_ sky130_fd_sc_hd__and2_1
XFILLER_119_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17298_ _01622_ _01623_ _01624_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__or3_1
XFILLER_174_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16249_ _08746_ _08747_ _08745_ vssd1 vssd1 vccd1 vccd1 _08861_ sky130_fd_sc_hd__a21bo_1
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19939_ net168 _00870_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18977__157 clknet_1_1__leaf__02729_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__inv_2
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10260_ _03191_ vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10191_ _03143_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__clkbuf_4
XFILLER_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13950_ _05380_ _06683_ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__or2_1
XFILLER_115_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12901_ _05508_ _05654_ _05655_ _05657_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__a22oi_2
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13881_ _05369_ _05333_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__nor2_4
XFILLER_189_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15620_ rbzero.debug_overlay.playerY\[-2\] rbzero.debug_overlay.playerX\[-2\] _06851_
+ vssd1 vssd1 vccd1 vccd1 _08304_ sky130_fd_sc_hd__mux2_1
X_12832_ _05492_ _05548_ _05553_ _05547_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__a22oi_2
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _07735_ _08108_ _08104_ _08103_ vssd1 vssd1 vccd1 vccd1 _08235_ sky130_fd_sc_hd__o31a_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _05505_ _05517_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__or2_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _07100_ _07123_ vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__nor2_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ net7 _04490_ _04491_ net6 vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__a31o_1
X_18270_ _02366_ vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__clkbuf_1
X_15482_ _08036_ _08038_ vssd1 vssd1 vccd1 vccd1 _08167_ sky130_fd_sc_hd__nor2_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _05309_ _05402_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__or2_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _01556_ _01557_ _01558_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__o21ai_1
X_14433_ _07119_ _07109_ _07120_ vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__or3_1
XFILLER_35_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11645_ _04424_ _04425_ _03739_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__mux2_1
XFILLER_161_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17152_ _09021_ _09046_ _09642_ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput15 i_gpout2_sel[0] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_8
X_14364_ _04840_ _06914_ _07032_ _07051_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__o31a_4
X_11576_ rbzero.tex_b0\[29\] rbzero.tex_b0\[28\] _03732_ vssd1 vssd1 vccd1 vccd1 _04358_
+ sky130_fd_sc_hd__mux2_1
Xinput26 i_gpout3_sel[5] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__buf_4
Xinput37 i_gpout5_sel[4] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_8
XFILLER_167_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput48 i_tex_in[1] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__buf_4
XFILLER_156_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16103_ _04946_ _08716_ vssd1 vssd1 vccd1 vccd1 _08717_ sky130_fd_sc_hd__nand2_1
X_13315_ _05472_ _06071_ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__nor2_1
X_17083_ _09660_ _09686_ vssd1 vssd1 vccd1 vccd1 _09688_ sky130_fd_sc_hd__or2_1
XFILLER_171_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__02741_ clknet_0__02741_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02741_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10527_ rbzero.tex_b0\[6\] rbzero.tex_b0\[5\] _03324_ vssd1 vssd1 vccd1 vccd1 _03331_
+ sky130_fd_sc_hd__mux2_1
X_14295_ rbzero.debug_overlay.playerY\[-3\] _06982_ _04928_ vssd1 vssd1 vccd1 vccd1
+ _06983_ sky130_fd_sc_hd__mux2_1
XFILLER_157_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16034_ _07494_ _07137_ _08647_ vssd1 vssd1 vccd1 vccd1 _08648_ sky130_fd_sc_hd__or3_1
X_10458_ rbzero.tex_b0\[39\] rbzero.tex_b0\[38\] _03291_ vssd1 vssd1 vccd1 vccd1 _03295_
+ sky130_fd_sc_hd__mux2_1
X_13246_ _05984_ _05985_ _05982_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__a21o_1
XFILLER_182_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10389_ rbzero.tex_b1\[7\] rbzero.tex_b1\[8\] _03254_ vssd1 vssd1 vccd1 vccd1 _03259_
+ sky130_fd_sc_hd__mux2_1
X_13177_ _05882_ _05933_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12128_ _04889_ _04862_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__xor2_1
X_17985_ _02193_ vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16936_ _09009_ _09007_ _09039_ _09035_ vssd1 vssd1 vccd1 vccd1 _09542_ sky130_fd_sc_hd__or4_1
X_19724_ clknet_leaf_95_i_clk _00655_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12059_ _04829_ vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16867_ _09472_ _09473_ vssd1 vssd1 vccd1 vccd1 _09474_ sky130_fd_sc_hd__nor2_1
X_19655_ clknet_leaf_17_i_clk _00586_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18606_ _02522_ vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__clkbuf_1
X_15818_ rbzero.traced_texa\[-1\] _08461_ _08459_ rbzero.wall_tracer.visualWallDist\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__a22o_1
X_19586_ clknet_leaf_61_i_clk _00517_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16798_ _09298_ _09299_ vssd1 vssd1 vccd1 vccd1 _09406_ sky130_fd_sc_hd__nor2_1
XFILLER_179_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18537_ _02486_ vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__clkbuf_1
X_15749_ rbzero.debug_overlay.playerY\[-1\] rbzero.debug_overlay.playerX\[-1\] _06851_
+ vssd1 vssd1 vccd1 vccd1 _08432_ sky130_fd_sc_hd__mux2_1
XFILLER_179_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18468_ _02450_ vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17419_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.wall_tracer.rayAddendY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__and2_1
XFILLER_53_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19178__338 clknet_1_1__leaf__02749_ vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__inv_2
XFILLER_14_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20430_ net490 _01361_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20361_ net421 _01292_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20292_ net352 _01223_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11430_ _03607_ _04209_ _04213_ _03627_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__a211o_1
XFILLER_137_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11361_ _03461_ _02904_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__nand2_1
XFILLER_193_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10312_ _03218_ vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__clkbuf_1
X_13100_ _05633_ _05639_ _05641_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__a21o_1
X_11292_ _04072_ _04073_ _04074_ _04076_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__a31o_1
X_14080_ rbzero.wall_tracer.trackDistX\[0\] _06788_ _06803_ vssd1 vssd1 vccd1 vccd1
+ _00439_ sky130_fd_sc_hd__o21a_1
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10243_ _03182_ vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__clkbuf_1
X_13031_ _05776_ _05786_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__or2b_1
XFILLER_152_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10174_ _03146_ vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17770_ _02014_ _02032_ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__or2b_1
X_14982_ _06787_ _07669_ vssd1 vssd1 vccd1 vccd1 _07670_ sky130_fd_sc_hd__nand2_1
XFILLER_121_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16721_ _09214_ _09219_ _09217_ vssd1 vssd1 vccd1 vccd1 _09329_ sky130_fd_sc_hd__a21oi_1
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13933_ _06675_ _05476_ _06684_ _06629_ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__a31o_1
XFILLER_47_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19440_ gpout2.clk_div\[0\] gpout2.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__or2_1
X_16652_ _09252_ _09260_ vssd1 vssd1 vccd1 vccd1 _09261_ sky130_fd_sc_hd__and2_1
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13864_ _06601_ _06620_ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__nor2_1
XFILLER_74_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15603_ _08115_ _08161_ _08159_ vssd1 vssd1 vccd1 vccd1 _08287_ sky130_fd_sc_hd__a21oi_2
XFILLER_90_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19371_ rbzero.traced_texa\[7\] rbzero.texV\[7\] vssd1 vssd1 vccd1 vccd1 _02850_
+ sky130_fd_sc_hd__nand2_1
X_12815_ _05510_ _05511_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__xnor2_1
X_16583_ _08844_ _09074_ _09192_ vssd1 vssd1 vccd1 vccd1 _09193_ sky130_fd_sc_hd__a21oi_1
XFILLER_15_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13795_ _06546_ _06547_ _06549_ _06551_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__a211o_1
XFILLER_16_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18322_ _02395_ vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__clkbuf_1
X_15534_ _08216_ _08217_ vssd1 vssd1 vccd1 vccd1 _08218_ sky130_fd_sc_hd__nor2_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12746_ _05502_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__clkbuf_4
XFILLER_188_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18253_ _04828_ vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__buf_4
XFILLER_163_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15465_ _08147_ _08148_ _08149_ vssd1 vssd1 vccd1 vccd1 _08150_ sky130_fd_sc_hd__or3_1
XFILLER_147_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12677_ _05314_ _05331_ _05315_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__mux2_1
X_17204_ _01541_ _01542_ _01543_ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__nand3_1
XFILLER_147_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14416_ _06733_ _07103_ vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__xnor2_1
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11628_ _03693_ _04408_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__or2_1
X_18184_ rbzero.spi_registers.got_new_leak _02262_ vssd1 vssd1 vccd1 vccd1 _02310_
+ sky130_fd_sc_hd__nand2_2
X_15396_ _07839_ vssd1 vssd1 vccd1 vccd1 _08081_ sky130_fd_sc_hd__clkbuf_4
XFILLER_200_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17135_ _09672_ _09685_ _01478_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__a21o_1
XFILLER_155_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14347_ _07034_ rbzero.debug_overlay.playerX\[-1\] _06887_ vssd1 vssd1 vccd1 vccd1
+ _07035_ sky130_fd_sc_hd__mux2_1
X_11559_ rbzero.tex_b0\[45\] rbzero.tex_b0\[44\] _04188_ vssd1 vssd1 vccd1 vccd1 _04341_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17066_ _08888_ _08317_ vssd1 vssd1 vccd1 vccd1 _09671_ sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1__f__02724_ clknet_0__02724_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02724_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14278_ _04947_ _06960_ _06964_ _06965_ vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_100_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16017_ _08629_ _08630_ vssd1 vssd1 vccd1 vccd1 _08631_ sky130_fd_sc_hd__nor2_1
Xclkbuf_0__02755_ _02755_ vssd1 vssd1 vccd1 vccd1 clknet_0__02755_ sky130_fd_sc_hd__clkbuf_16
XFILLER_131_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13229_ _05984_ _05985_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__xor2_4
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17968_ _02184_ vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19707_ clknet_leaf_71_i_clk _00638_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16919_ _08512_ _09525_ _08489_ vssd1 vssd1 vccd1 vccd1 _09526_ sky130_fd_sc_hd__a21oi_1
XFILLER_65_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17899_ _02148_ vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19638_ clknet_leaf_38_i_clk _00569_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19569_ clknet_leaf_36_i_clk _00500_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20413_ net473 _01344_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20344_ net404 _01275_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20275_ net335 _01206_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10930_ _03583_ _03582_ _03598_ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__o21a_1
XFILLER_5_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__02744_ clknet_0__02744_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02744_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_147_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10861_ _03619_ _03633_ _03646_ _03540_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__a211o_1
XFILLER_147_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ _05253_ _05257_ _05311_ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__mux2_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _05527_ _05992_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__nor2_1
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10792_ rbzero.traced_texVinit\[7\] rbzero.spi_registers.vshift\[4\] vssd1 vssd1
+ vccd1 vccd1 _03578_ sky130_fd_sc_hd__or2_1
XFILLER_25_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _05178_ _05180_ _05181_ _05174_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__a31o_1
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15250_ _07936_ _04923_ _06851_ vssd1 vssd1 vccd1 vccd1 _07937_ sky130_fd_sc_hd__mux2_2
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12462_ _05131_ _05218_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__xnor2_4
XFILLER_12_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14201_ rbzero.debug_overlay.playerX\[-8\] rbzero.debug_overlay.playerX\[-9\] rbzero.debug_overlay.playerX\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__o21ai_1
X_11413_ _03671_ _04191_ _04196_ _03648_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__a211o_1
XFILLER_172_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_82 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_82/HI o_rgb[11] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_93 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_93/HI zeros[2] sky130_fd_sc_hd__conb_1
XFILLER_172_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15181_ _07864_ _07866_ vssd1 vssd1 vccd1 vccd1 _07868_ sky130_fd_sc_hd__nand2_1
XFILLER_32_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12393_ _05081_ _05133_ _05147_ _05149_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__nor4b_2
XFILLER_137_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14132_ rbzero.wall_tracer.stepDistX\[3\] _06753_ _06825_ vssd1 vssd1 vccd1 vccd1
+ _06831_ sky130_fd_sc_hd__mux2_1
XFILLER_181_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11344_ rbzero.debug_overlay.playerX\[2\] _04068_ _04092_ rbzero.debug_overlay.playerX\[-3\]
+ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__a22o_1
XFILLER_67_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14063_ rbzero.wall_tracer.visualWallDist\[-7\] _03496_ _06791_ rbzero.wall_tracer.trackDistX\[-7\]
+ _03485_ vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__o221a_1
X_11275_ _04052_ _04054_ _04040_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__nand3b_2
XFILLER_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13014_ _05516_ _05610_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__nor2_1
X_10226_ _03173_ vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__02440_ clknet_0__02440_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02440_
+ sky130_fd_sc_hd__clkbuf_16
X_18871_ rbzero.hsync _02700_ _02701_ vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__o21a_1
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10157_ rbzero.tex_g0\[54\] rbzero.tex_g0\[53\] _03132_ vssd1 vssd1 vccd1 vccd1 _03137_
+ sky130_fd_sc_hd__mux2_1
X_17822_ _02073_ _02074_ _02084_ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__nand3_1
XFILLER_94_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10088_ rbzero.tex_g1\[22\] rbzero.tex_g1\[23\] _03095_ vssd1 vssd1 vccd1 vccd1 _03101_
+ sky130_fd_sc_hd__mux2_1
X_14965_ _07623_ _07652_ vssd1 vssd1 vccd1 vccd1 _07653_ sky130_fd_sc_hd__xor2_1
X_17753_ _02005_ _02006_ _02021_ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__a21o_1
X_13916_ rbzero.wall_tracer.stepDistY\[-8\] _06669_ _00004_ vssd1 vssd1 vccd1 vccd1
+ _06670_ sky130_fd_sc_hd__mux2_1
X_16704_ _09309_ _09310_ _09311_ vssd1 vssd1 vccd1 vccd1 _09313_ sky130_fd_sc_hd__o21ai_1
X_17684_ rbzero.debug_overlay.vplaneX\[-6\] _01948_ vssd1 vssd1 vccd1 vccd1 _01958_
+ sky130_fd_sc_hd__nand2_1
XFILLER_35_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14896_ _07550_ _07561_ vssd1 vssd1 vccd1 vccd1 _07584_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16635_ _09213_ _09243_ vssd1 vssd1 vccd1 vccd1 _09244_ sky130_fd_sc_hd__xnor2_1
X_19423_ _08452_ _01921_ _02880_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__and3_1
XFILLER_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13847_ _06589_ _06602_ _06603_ vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__mux2_1
X_16566_ _09058_ _09059_ vssd1 vssd1 vccd1 vccd1 _09176_ sky130_fd_sc_hd__and2b_1
X_19354_ _02829_ _02832_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__nand2_1
XFILLER_188_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13778_ _06521_ _06534_ vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__nand2_1
XFILLER_149_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15517_ _08199_ _08200_ vssd1 vssd1 vccd1 vccd1 _08201_ sky130_fd_sc_hd__and2_1
X_18305_ _02379_ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__inv_2
X_12729_ _05481_ _05485_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__xnor2_1
X_19285_ rbzero.traced_texa\[-7\] rbzero.texV\[-7\] vssd1 vssd1 vccd1 vccd1 _02778_
+ sky130_fd_sc_hd__and2_1
X_16497_ _09105_ _09106_ vssd1 vssd1 vccd1 vccd1 _09107_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18236_ _02345_ vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__clkbuf_1
X_15448_ _07756_ vssd1 vssd1 vccd1 vccd1 _08133_ sky130_fd_sc_hd__buf_2
XFILLER_31_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18167_ rbzero.spi_registers.new_mapd\[5\] _02290_ _02300_ _02301_ vssd1 vssd1 vccd1
+ vccd1 _00768_ sky130_fd_sc_hd__o211a_1
X_15379_ _08045_ _08046_ vssd1 vssd1 vccd1 vccd1 _08064_ sky130_fd_sc_hd__or2_1
XFILLER_129_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17118_ _09649_ vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__inv_2
X_18098_ net44 rbzero.spi_registers.sclk_buffer\[0\] _03337_ vssd1 vssd1 vccd1 vccd1
+ _02254_ sky130_fd_sc_hd__mux2_1
XFILLER_172_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09940_ rbzero.tex_r0\[29\] rbzero.tex_r0\[28\] _03017_ vssd1 vssd1 vccd1 vccd1 _03023_
+ sky130_fd_sc_hd__mux2_1
X_17049_ _09280_ _09634_ _09653_ vssd1 vssd1 vccd1 vccd1 _09654_ sky130_fd_sc_hd__o21ai_1
XFILLER_171_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__02738_ _02738_ vssd1 vssd1 vccd1 vccd1 clknet_0__02738_ sky130_fd_sc_hd__clkbuf_16
X_20060_ clknet_leaf_1_i_clk _00991_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ss_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_09871_ rbzero.tex_r0\[62\] rbzero.tex_r0\[61\] _02984_ vssd1 vssd1 vccd1 vccd1 _02987_
+ sky130_fd_sc_hd__mux2_1
XFILLER_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20327_ net387 _01258_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11060_ rbzero.debug_overlay.playerX\[0\] _03462_ _03474_ rbzero.debug_overlay.playerX\[3\]
+ _03845_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__a221o_1
X_20258_ net318 _01189_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10011_ rbzero.tex_g1\[58\] rbzero.tex_g1\[59\] _02976_ vssd1 vssd1 vccd1 vccd1 _03060_
+ sky130_fd_sc_hd__mux2_1
XFILLER_135_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20189_ net249 _01120_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_49_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ _07434_ _07437_ _07436_ vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__a21oi_1
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11962_ net29 _04729_ _04735_ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__a21oi_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _06452_ _06457_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__or2b_1
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10913_ _03614_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__buf_6
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ _07339_ _07368_ vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__nor2_1
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ net21 net22 vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__and2b_1
XFILLER_189_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__02727_ clknet_0__02727_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02727_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_72_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16420_ _08913_ _08915_ _08912_ vssd1 vssd1 vccd1 vccd1 _09031_ sky130_fd_sc_hd__a21bo_1
X_13632_ _06125_ _06383_ _06388_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__a21oi_1
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10844_ _03626_ _03629_ rbzero.row_render.texu\[0\] vssd1 vssd1 vccd1 vccd1 _03630_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_73_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16351_ _08960_ _08961_ _08962_ vssd1 vssd1 vccd1 vccd1 _08963_ sky130_fd_sc_hd__a21o_1
X_13563_ _06312_ _06318_ _06319_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__a21boi_1
X_10775_ _03559_ _03560_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__nor2_1
XFILLER_73_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15302_ _07978_ _07986_ vssd1 vssd1 vccd1 vccd1 _07988_ sky130_fd_sc_hd__or2_1
XFILLER_9_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12514_ _05270_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__buf_2
X_16282_ _08893_ vssd1 vssd1 vccd1 vccd1 _08894_ sky130_fd_sc_hd__clkinv_2
XFILLER_158_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13494_ _06244_ _06249_ _06250_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__o21a_1
XFILLER_160_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18021_ _02212_ vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__clkbuf_1
X_15233_ _07780_ _07798_ _07778_ vssd1 vssd1 vccd1 vccd1 _07920_ sky130_fd_sc_hd__a21oi_1
XFILLER_201_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12445_ _05077_ _05195_ _05149_ _05153_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__a211o_1
XFILLER_60_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15164_ _07712_ _07722_ _07720_ vssd1 vssd1 vccd1 vccd1 _07851_ sky130_fd_sc_hd__a21o_1
XFILLER_126_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12376_ _05087_ _05089_ _05094_ _05132_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__a211o_2
XFILLER_114_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14115_ rbzero.wall_tracer.stepDistX\[-5\] _06695_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _06822_ sky130_fd_sc_hd__mux2_1
XFILLER_141_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11327_ rbzero.debug_overlay.vplaneY\[-1\] _04093_ _04056_ _04109_ _04111_ vssd1
+ vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__a221o_1
X_19972_ net201 _00903_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[52\] sky130_fd_sc_hd__dfxtp_1
X_15095_ _07267_ _07271_ _07264_ vssd1 vssd1 vccd1 vccd1 _07783_ sky130_fd_sc_hd__a21bo_1
XFILLER_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14046_ rbzero.wall_tracer.stepDistY\[10\] _06781_ _04836_ vssd1 vssd1 vccd1 vccd1
+ _06782_ sky130_fd_sc_hd__mux2_1
XFILLER_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11258_ _03512_ _04042_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__nor2_1
X_19236__11 clknet_1_1__leaf__02754_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__inv_2
X_10209_ _03164_ vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18854_ rbzero.pov.ready_buffer\[8\] _02635_ _02689_ _02672_ vssd1 vssd1 vccd1 vccd1
+ _01067_ sky130_fd_sc_hd__o211a_1
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11189_ rbzero.tex_r1\[9\] _03919_ _03926_ _03670_ vssd1 vssd1 vccd1 vccd1 _03974_
+ sky130_fd_sc_hd__a31o_1
XFILLER_121_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17805_ _02000_ rbzero.debug_overlay.vplaneX\[-1\] vssd1 vssd1 vccd1 vccd1 _02070_
+ sky130_fd_sc_hd__nor2_1
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15997_ _08607_ _08610_ vssd1 vssd1 vccd1 vccd1 _08611_ sky130_fd_sc_hd__xnor2_1
X_18785_ rbzero.pov.ready_buffer\[42\] _02636_ _02652_ _02643_ vssd1 vssd1 vccd1 vccd1
+ _01035_ sky130_fd_sc_hd__o211a_1
XFILLER_83_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19251__25 clknet_1_1__leaf__02755_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__inv_2
XFILLER_83_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14948_ _07614_ _07635_ vssd1 vssd1 vccd1 vccd1 _07636_ sky130_fd_sc_hd__or2_1
X_17736_ _01977_ _01992_ _01993_ _01997_ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__o31ai_1
XFILLER_91_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14879_ _07547_ _07566_ _07564_ vssd1 vssd1 vccd1 vccd1 _07567_ sky130_fd_sc_hd__a21o_1
X_17667_ rbzero.debug_overlay.vplaneX\[-3\] rbzero.wall_tracer.rayAddendX\[-3\] vssd1
+ vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__nor2_1
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19406_ gpout0.clk_div\[0\] gpout0.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__nand2_1
X_16618_ _09114_ _09116_ _09113_ vssd1 vssd1 vccd1 vccd1 _09227_ sky130_fd_sc_hd__a21bo_1
XFILLER_126_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17598_ rbzero.wall_tracer.rayAddendY\[8\] rbzero.wall_tracer.rayAddendY\[7\] _01785_
+ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__o21ai_1
XFILLER_50_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16549_ _07992_ _09035_ vssd1 vssd1 vccd1 vccd1 _09159_ sky130_fd_sc_hd__nor2_1
X_19337_ _02759_ _02820_ _02821_ _02319_ rbzero.texV\[1\] vssd1 vssd1 vccd1 vccd1
+ _01418_ sky130_fd_sc_hd__a32o_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19268_ rbzero.traced_texa\[-10\] rbzero.texV\[-10\] vssd1 vssd1 vccd1 vccd1 _02764_
+ sky130_fd_sc_hd__nand2_1
XFILLER_148_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18219_ _02333_ vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20112_ clknet_leaf_90_i_clk _01043_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
X_09923_ rbzero.tex_r0\[37\] rbzero.tex_r0\[36\] _03006_ vssd1 vssd1 vccd1 vccd1 _03014_
+ sky130_fd_sc_hd__mux2_1
XFILLER_131_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20043_ clknet_leaf_7_i_clk _00974_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_09854_ _02909_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__clkbuf_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09785_ rbzero.tex_r1\[36\] rbzero.tex_r1\[37\] _02932_ vssd1 vssd1 vccd1 vccd1 _02940_
+ sky130_fd_sc_hd__mux2_1
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18435__75 clknet_1_1__leaf__02438_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__inv_2
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10560_ _03350_ rbzero.map_rom.i_col\[4\] _03351_ rbzero.debug_overlay.playerY\[5\]
+ _03355_ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__a221o_1
XFILLER_167_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10491_ rbzero.tex_b0\[23\] rbzero.tex_b0\[22\] _03302_ vssd1 vssd1 vccd1 vccd1 _03312_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12230_ _04969_ _04987_ _04988_ _04967_ _04965_ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__a32o_1
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12161_ _04922_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_31_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_107_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11112_ _03848_ _03887_ _03897_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__a21o_1
XFILLER_107_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12092_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__nand2_1
XFILLER_151_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11043_ rbzero.floor_leak\[5\] _03718_ _03828_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__a21oi_1
XFILLER_122_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15920_ rbzero.wall_tracer.trackDistX\[-7\] rbzero.wall_tracer.stepDistX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _08541_ sky130_fd_sc_hd__and2_1
XFILLER_104_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_46_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_15851_ _08468_ _08471_ _08480_ vssd1 vssd1 vccd1 vccd1 _08481_ sky130_fd_sc_hd__and3_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _06871_ _06966_ _07048_ _06949_ vssd1 vssd1 vccd1 vccd1 _07490_ sky130_fd_sc_hd__o22ai_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18570_ rbzero.pov.spi_buffer\[53\] rbzero.pov.spi_buffer\[54\] _02499_ vssd1 vssd1
+ vccd1 vccd1 _02504_ sky130_fd_sc_hd__mux2_1
X_15782_ rbzero.row_render.side _08449_ _08453_ _06851_ vssd1 vssd1 vccd1 vccd1 _00491_
+ sky130_fd_sc_hd__a22o_1
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12994_ _05713_ _05714_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17521_ _01803_ _01810_ _01804_ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__nand3_1
X_14733_ _07419_ _07420_ vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__nor2_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11945_ net25 net26 _04719_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__and3b_1
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__nand2_1
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14664_ _06921_ _07351_ vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__xnor2_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ _04503_ _03902_ _04612_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__mux2_1
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16403_ _07494_ vssd1 vssd1 vccd1 vccd1 _09014_ sky130_fd_sc_hd__buf_2
XFILLER_177_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13615_ _06364_ _06365_ _06371_ vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__a21o_1
X_10827_ _03552_ _03555_ _03603_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__a21oi_2
X_17383_ _08474_ _08477_ vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__xor2_1
X_14595_ _07280_ _07282_ vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__nor2_1
XFILLER_164_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16334_ _08943_ _08945_ vssd1 vssd1 vccd1 vccd1 _08946_ sky130_fd_sc_hd__xor2_1
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13546_ _06232_ _06234_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__xnor2_1
X_10758_ rbzero.texV\[4\] _03542_ _03543_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__nand3_1
XFILLER_119_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16265_ _08875_ _08876_ vssd1 vssd1 vccd1 vccd1 _08877_ sky130_fd_sc_hd__nor2_1
XFILLER_125_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13477_ _06158_ _06233_ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__and2_1
X_10689_ rbzero.wall_tracer.state\[8\] vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__inv_2
XFILLER_127_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15216_ _07892_ _07902_ vssd1 vssd1 vccd1 vccd1 _07903_ sky130_fd_sc_hd__xnor2_1
X_18004_ _02203_ vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12428_ _05158_ _05175_ _05182_ _05184_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__and4b_1
XFILLER_161_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16196_ _08679_ _08685_ vssd1 vssd1 vccd1 vccd1 _08809_ sky130_fd_sc_hd__nor2_1
XFILLER_160_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15147_ _07265_ _07270_ _07710_ vssd1 vssd1 vccd1 vccd1 _07834_ sky130_fd_sc_hd__or3_1
XFILLER_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12359_ rbzero.wall_tracer.rayAddendX\[-3\] _05115_ _05072_ vssd1 vssd1 vccd1 vccd1
+ _05116_ sky130_fd_sc_hd__mux2_2
XFILLER_114_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19955_ net184 _00886_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[35\] sky130_fd_sc_hd__dfxtp_1
X_15078_ _07198_ vssd1 vssd1 vccd1 vccd1 _07766_ sky130_fd_sc_hd__clkbuf_4
XFILLER_45_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14029_ _06768_ vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19886_ clknet_leaf_23_i_clk _00817_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_67_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18837_ _01752_ _02635_ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__nand2_1
XFILLER_68_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__02437_ _02437_ vssd1 vssd1 vccd1 vccd1 clknet_0__02437_ sky130_fd_sc_hd__clkbuf_16
XFILLER_55_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18768_ rbzero.debug_overlay.facingX\[-6\] _02638_ vssd1 vssd1 vccd1 vccd1 _02642_
+ sky130_fd_sc_hd__or2_1
XFILLER_67_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17719_ _01974_ _01988_ _01987_ _01986_ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__o211ai_2
X_18699_ _02589_ _06909_ _02539_ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__mux2_1
XFILLER_50_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09906_ rbzero.tex_r0\[45\] rbzero.tex_r0\[44\] _02995_ vssd1 vssd1 vccd1 vccd1 _03005_
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20026_ clknet_leaf_86_i_clk _00957_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_09837_ _02967_ vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09768_ rbzero.tex_r1\[44\] rbzero.tex_r1\[45\] _02921_ vssd1 vssd1 vccd1 vccd1 _02931_
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _03517_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__clkbuf_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11661_ rbzero.tex_b1\[17\] rbzero.tex_b1\[16\] _04376_ vssd1 vssd1 vccd1 vccd1 _04442_
+ sky130_fd_sc_hd__mux2_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13400_ _05990_ _06156_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__nor2_1
X_10612_ _03398_ _03405_ _03407_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__nand3b_1
X_14380_ _06871_ _07024_ _07037_ _07047_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__or4_1
X_11592_ rbzero.tex_b0\[7\] rbzero.tex_b0\[6\] _03699_ vssd1 vssd1 vccd1 vccd1 _04374_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13331_ _06008_ _06061_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__nor2_1
XFILLER_155_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10543_ net72 _02907_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__nand2_4
XFILLER_183_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16050_ _07530_ _08133_ _08380_ vssd1 vssd1 vccd1 vccd1 _08664_ sky130_fd_sc_hd__o21ai_1
XFILLER_155_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13262_ _05965_ _06018_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__xor2_1
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10474_ _03303_ vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__clkbuf_1
XFILLER_157_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15001_ _07612_ _07638_ _07643_ _07688_ vssd1 vssd1 vccd1 vccd1 _07689_ sky130_fd_sc_hd__and4_1
X_12213_ rbzero.wall_tracer.trackDistY\[-9\] vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__inv_2
XFILLER_142_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13193_ _05906_ _05949_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__or2_2
XFILLER_159_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12144_ _04899_ _04853_ _04867_ _04848_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__o211ai_1
XFILLER_111_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19740_ clknet_leaf_76_i_clk _00671_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_16952_ _09545_ _09557_ vssd1 vssd1 vccd1 vccd1 _09558_ sky130_fd_sc_hd__xor2_1
XFILLER_150_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12075_ _04838_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__clkbuf_4
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11026_ rbzero.row_render.size\[2\] gpout0.hpos\[2\] _03501_ _03811_ vssd1 vssd1
+ vccd1 vccd1 _03812_ sky130_fd_sc_hd__a211o_1
X_15903_ _08519_ _08520_ vssd1 vssd1 vccd1 vccd1 _08526_ sky130_fd_sc_hd__and2_1
X_19671_ clknet_leaf_34_i_clk _00602_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.i_col\[4\]
+ sky130_fd_sc_hd__dfxtp_4
X_16883_ _09488_ _09489_ vssd1 vssd1 vccd1 vccd1 _09490_ sky130_fd_sc_hd__xnor2_2
XFILLER_37_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18622_ _02530_ vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__clkbuf_1
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15834_ _08465_ vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__clkbuf_1
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18414__56 clknet_1_1__leaf__02436_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__inv_2
XFILLER_92_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18553_ rbzero.pov.spi_buffer\[45\] rbzero.pov.spi_buffer\[46\] _02488_ vssd1 vssd1
+ vccd1 vccd1 _02495_ sky130_fd_sc_hd__mux2_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12977_ _05704_ _05706_ _05705_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__a21o_1
X_15765_ net61 _04054_ vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__nor2_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ _01714_ _01795_ _08448_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__a21o_1
XFILLER_166_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14716_ _07395_ _07399_ _07403_ vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__a21o_1
X_11928_ net25 _04701_ _04702_ net24 vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__a31o_1
X_15696_ _08261_ _08263_ _08259_ vssd1 vssd1 vccd1 vccd1 _08379_ sky130_fd_sc_hd__a21bo_1
X_18484_ rbzero.pov.spi_buffer\[12\] rbzero.pov.spi_buffer\[13\] _02455_ vssd1 vssd1
+ vccd1 vccd1 _02459_ sky130_fd_sc_hd__mux2_1
XFILLER_178_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14647_ _07331_ _07334_ vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__xnor2_2
X_17435_ rbzero.debug_overlay.vplaneY\[-7\] _01723_ vssd1 vssd1 vccd1 vccd1 _01732_
+ sky130_fd_sc_hd__or2_1
X_11859_ net12 _04624_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__nor2_2
XFILLER_60_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_18 rbzero.debug_overlay.facingX\[-1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14578_ _06857_ _07007_ vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__nor2_1
XANTENNA_29 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17366_ _01675_ vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__clkbuf_1
X_16317_ _08927_ _08928_ vssd1 vssd1 vccd1 vccd1 _08929_ sky130_fd_sc_hd__nor2_1
XFILLER_159_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13529_ _06275_ _06273_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__xor2_1
XFILLER_158_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17297_ _01617_ _01619_ _01616_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__a21boi_2
X_16248_ _08858_ _08859_ vssd1 vssd1 vccd1 vccd1 _08860_ sky130_fd_sc_hd__xor2_1
XFILLER_174_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16179_ _07992_ _08133_ vssd1 vssd1 vccd1 vccd1 _08792_ sky130_fd_sc_hd__nor2_1
XFILLER_161_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19938_ net167 _00869_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19869_ clknet_leaf_20_i_clk _00800_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19155__317 clknet_1_1__leaf__02747_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__inv_2
XFILLER_137_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10190_ _03154_ vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12900_ _05504_ _05656_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__xnor2_1
X_20009_ clknet_leaf_75_i_clk _00940_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_19049__222 clknet_1_1__leaf__02736_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__inv_2
X_13880_ _06633_ _06635_ _06603_ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__mux2_1
XFILLER_101_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12831_ _05475_ _05486_ _05587_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__a21o_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15550_ _08232_ _08233_ vssd1 vssd1 vccd1 vccd1 _08234_ sky130_fd_sc_hd__xnor2_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _05513_ _05518_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__or2_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _07143_ _07188_ vssd1 vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__xnor2_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _04487_ net62 vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__or2_1
X_15481_ _08093_ _08165_ vssd1 vssd1 vccd1 vccd1 _08166_ sky130_fd_sc_hd__xnor2_2
XFILLER_70_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12693_ _05404_ _05425_ _05433_ _05443_ _05449_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__a2111o_4
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _01522_ vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__clkbuf_4
X_14432_ _07101_ _07117_ vssd1 vssd1 vccd1 vccd1 _07120_ sky130_fd_sc_hd__or2_1
XFILLER_175_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11644_ rbzero.tex_b1\[51\] rbzero.tex_b1\[50\] _04376_ vssd1 vssd1 vccd1 vccd1 _04425_
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17151_ _09674_ _09679_ _09681_ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__a21oi_1
XFILLER_126_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14363_ rbzero.wall_tracer.visualWallDist\[0\] _06855_ _07050_ _04948_ vssd1 vssd1
+ vccd1 vccd1 _07051_ sky130_fd_sc_hd__o2bb2a_1
X_11575_ _04198_ _04352_ _04356_ _03704_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__a211o_1
XFILLER_7_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput16 i_gpout2_sel[1] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_6
Xinput27 i_gpout4_sel[0] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_4
XFILLER_35_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16102_ _08713_ _08715_ vssd1 vssd1 vccd1 vccd1 _08716_ sky130_fd_sc_hd__xor2_2
XFILLER_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput38 i_gpout5_sel[5] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_4
X_13314_ _06070_ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__clkbuf_4
Xinput49 i_tex_in[2] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_6
X_17082_ _09660_ _09686_ vssd1 vssd1 vccd1 vccd1 _09687_ sky130_fd_sc_hd__nand2_1
X_10526_ _03330_ vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__02740_ clknet_0__02740_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02740_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_182_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19095__264 clknet_1_1__leaf__02740_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__inv_2
XFILLER_128_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14294_ _06980_ _06981_ vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__and2_1
XFILLER_183_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16033_ _07273_ _07198_ vssd1 vssd1 vccd1 vccd1 _08647_ sky130_fd_sc_hd__or2_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13245_ _05950_ _05986_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__nor2_4
XFILLER_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10457_ _03294_ vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__clkbuf_1
X_13176_ _05925_ _05932_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__xor2_1
X_10388_ _03258_ vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12127_ _04863_ _04858_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__and2b_1
X_17984_ rbzero.pov.spi_buffer\[45\] rbzero.pov.ready_buffer\[45\] _02186_ vssd1 vssd1
+ vccd1 vccd1 _02193_ sky130_fd_sc_hd__mux2_1
XFILLER_81_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19723_ clknet_leaf_87_i_clk _00654_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16935_ _09009_ _09035_ vssd1 vssd1 vccd1 vccd1 _09541_ sky130_fd_sc_hd__nor2_1
X_12058_ net72 rbzero.wall_tracer.state\[2\] _04828_ vssd1 vssd1 vccd1 vccd1 _04829_
+ sky130_fd_sc_hd__and3_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11009_ _02902_ _03780_ _03793_ gpout0.hpos\[9\] _03794_ vssd1 vssd1 vccd1 vccd1
+ _03795_ sky130_fd_sc_hd__o221a_1
X_19654_ clknet_leaf_18_i_clk _00585_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16866_ _09283_ _09385_ _09280_ vssd1 vssd1 vccd1 vccd1 _09473_ sky130_fd_sc_hd__a21boi_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18605_ rbzero.pov.spi_buffer\[70\] rbzero.pov.spi_buffer\[71\] _02443_ vssd1 vssd1
+ vccd1 vccd1 _02522_ sky130_fd_sc_hd__mux2_1
X_15817_ rbzero.traced_texa\[-2\] _08461_ _08459_ rbzero.wall_tracer.visualWallDist\[-2\]
+ vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__a22o_1
XFILLER_19_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19585_ clknet_leaf_61_i_clk _00516_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16797_ _09403_ _09404_ vssd1 vssd1 vccd1 vccd1 _09405_ sky130_fd_sc_hd__nand2_1
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18536_ rbzero.pov.spi_buffer\[37\] rbzero.pov.spi_buffer\[38\] _02477_ vssd1 vssd1
+ vccd1 vccd1 _02486_ sky130_fd_sc_hd__mux2_1
XFILLER_52_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15748_ _08312_ _08430_ vssd1 vssd1 vccd1 vccd1 _08431_ sky130_fd_sc_hd__xor2_4
XFILLER_52_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18467_ rbzero.pov.spi_buffer\[4\] rbzero.pov.spi_buffer\[5\] _02444_ vssd1 vssd1
+ vccd1 vccd1 _02450_ sky130_fd_sc_hd__mux2_1
X_15679_ _08224_ _08361_ vssd1 vssd1 vccd1 vccd1 _08362_ sky130_fd_sc_hd__nand2_1
XFILLER_21_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17418_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.wall_tracer.rayAddendY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__nor2_1
XFILLER_178_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17349_ rbzero.spi_registers.new_mapd\[3\] rbzero.spi_registers.spi_buffer\[3\] _01663_
+ vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__mux2_1
XFILLER_53_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20360_ net420 _01291_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20291_ net351 _01222_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11360_ _03519_ _04124_ _04144_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__a21bo_1
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10311_ rbzero.tex_b1\[44\] rbzero.tex_b1\[45\] _03210_ vssd1 vssd1 vccd1 vccd1 _03218_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11291_ _04037_ _04075_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__xnor2_2
XFILLER_106_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20489_ clknet_leaf_42_i_clk _01420_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13030_ _05776_ _05786_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10242_ rbzero.tex_g0\[14\] rbzero.tex_g0\[13\] _03177_ vssd1 vssd1 vccd1 vccd1 _03182_
+ sky130_fd_sc_hd__mux2_1
XFILLER_191_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10173_ rbzero.tex_g0\[47\] rbzero.tex_g0\[46\] _03144_ vssd1 vssd1 vccd1 vccd1 _03146_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14981_ _06872_ _07199_ vssd1 vssd1 vccd1 vccd1 _07669_ sky130_fd_sc_hd__nor2_1
XFILLER_102_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16720_ _09324_ _09327_ vssd1 vssd1 vccd1 vccd1 _09328_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13932_ _06665_ _06683_ _06664_ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__mux2_1
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16651_ _09258_ _09259_ vssd1 vssd1 vccd1 vccd1 _09260_ sky130_fd_sc_hd__xor2_1
X_13863_ _06573_ _06568_ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15602_ _08284_ _08285_ vssd1 vssd1 vccd1 vccd1 _08286_ sky130_fd_sc_hd__nand2_1
X_12814_ _05555_ _05570_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__xnor2_1
X_19370_ rbzero.traced_texa\[7\] rbzero.texV\[7\] vssd1 vssd1 vccd1 vccd1 _02849_
+ sky130_fd_sc_hd__nor2_1
X_16582_ _09071_ _09073_ vssd1 vssd1 vccd1 vccd1 _09192_ sky130_fd_sc_hd__nor2_1
X_13794_ _06537_ _06550_ vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__nand2_1
XFILLER_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18321_ rbzero.spi_registers.new_other\[7\] rbzero.spi_registers.spi_buffer\[7\]
+ _02388_ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__mux2_1
X_15533_ _08214_ _08215_ vssd1 vssd1 vccd1 vccd1 _08217_ sky130_fd_sc_hd__and2_1
X_12745_ _05450_ _05458_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__xnor2_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15464_ _07900_ _08019_ _08021_ _08012_ vssd1 vssd1 vccd1 vccd1 _08149_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18252_ rbzero.spi_registers.vshift\[5\] _02349_ vssd1 vssd1 vccd1 vccd1 _02355_
+ sky130_fd_sc_hd__or2_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12676_ _05209_ _05430_ _05431_ _05323_ _05432_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__a32oi_4
XFILLER_124_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17203_ _01535_ _01536_ _01537_ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__o21bai_1
X_14415_ _05414_ _06720_ _06725_ _06717_ vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__a211o_2
X_11627_ rbzero.tex_b1\[37\] rbzero.tex_b1\[36\] _03616_ vssd1 vssd1 vccd1 vccd1 _04408_
+ sky130_fd_sc_hd__mux2_1
X_19103__271 clknet_1_0__leaf__02741_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__inv_2
X_15395_ _08077_ _08078_ _08079_ vssd1 vssd1 vccd1 vccd1 _08080_ sky130_fd_sc_hd__o21a_1
X_18183_ rbzero.spi_registers.new_mapd\[1\] _02289_ _02309_ _02301_ vssd1 vssd1 vccd1
+ vccd1 _00776_ sky130_fd_sc_hd__o211a_1
XFILLER_200_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17134_ _09683_ _09684_ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__and2b_1
X_14346_ _07032_ _07033_ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__and2_1
X_11558_ rbzero.tex_b0\[47\] rbzero.tex_b0\[46\] _03699_ vssd1 vssd1 vccd1 vccd1 _04340_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17065_ _09668_ _09669_ vssd1 vssd1 vccd1 vccd1 _09670_ sky130_fd_sc_hd__nor2_1
X_10509_ _03321_ vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__02723_ clknet_0__02723_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02723_
+ sky130_fd_sc_hd__clkbuf_16
X_14277_ rbzero.debug_overlay.playerX\[-4\] _06887_ _04838_ vssd1 vssd1 vccd1 vccd1
+ _06965_ sky130_fd_sc_hd__a21oi_1
XFILLER_109_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11489_ _03671_ _04267_ _04271_ _03648_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__a211o_1
X_16016_ _08627_ _08628_ vssd1 vssd1 vccd1 vccd1 _08630_ sky130_fd_sc_hd__and2_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__02754_ _02754_ vssd1 vssd1 vccd1 vccd1 clknet_0__02754_ sky130_fd_sc_hd__clkbuf_16
X_13228_ _05944_ _05946_ _05948_ _05907_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__a22o_2
XFILLER_170_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13159_ _05914_ _05915_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__xnor2_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ rbzero.pov.spi_buffer\[37\] rbzero.pov.ready_buffer\[37\] _02175_ vssd1 vssd1
+ vccd1 vccd1 _02184_ sky130_fd_sc_hd__mux2_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19706_ clknet_leaf_71_i_clk _00637_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_16918_ _09523_ _09524_ vssd1 vssd1 vccd1 vccd1 _09525_ sky130_fd_sc_hd__xnor2_1
XFILLER_78_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17898_ rbzero.pov.spi_buffer\[4\] rbzero.pov.ready_buffer\[4\] _02143_ vssd1 vssd1
+ vccd1 vccd1 _02148_ sky130_fd_sc_hd__mux2_1
XFILLER_38_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19637_ clknet_leaf_38_i_clk _00568_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16849_ _09454_ _09455_ vssd1 vssd1 vccd1 vccd1 _09456_ sky130_fd_sc_hd__nor2_1
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19568_ clknet_leaf_36_i_clk _00499_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18519_ _02443_ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__clkbuf_4
XFILLER_178_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19499_ clknet_leaf_46_i_clk _00445_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[6\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20412_ net472 _01343_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20343_ net403 _01274_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20274_ net334 _01205_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__02743_ clknet_0__02743_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02743_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_186_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10860_ _03632_ _03645_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__nor2_1
XFILLER_71_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10791_ rbzero.traced_texVinit\[7\] rbzero.spi_registers.vshift\[4\] vssd1 vssd1
+ vccd1 vccd1 _03577_ sky130_fd_sc_hd__nand2_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _05221_ _05222_ _05223_ _05254_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__nor4_1
XFILLER_200_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ _05105_ _05127_ _05199_ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__o21a_1
XFILLER_200_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14200_ rbzero.debug_overlay.playerX\[-7\] rbzero.debug_overlay.playerX\[-8\] rbzero.debug_overlay.playerX\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__or3_1
X_11412_ _04192_ _04193_ _04194_ _04195_ _03607_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__o221a_1
XFILLER_149_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15180_ _07864_ _07866_ vssd1 vssd1 vccd1 vccd1 _07867_ sky130_fd_sc_hd__nor2_1
XFILLER_137_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtop_ew_algofoogle_83 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_83/HI o_rgb[12] sky130_fd_sc_hd__conb_1
X_12392_ _03488_ _05078_ _05148_ _05080_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__o31a_1
Xtop_ew_algofoogle_94 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_94/HI zeros[3] sky130_fd_sc_hd__conb_1
XFILLER_193_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14131_ _06830_ vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_193_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11343_ rbzero.debug_overlay.playerX\[-1\] _04093_ _04084_ rbzero.debug_overlay.playerX\[-6\]
+ _04127_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__a221o_1
XFILLER_192_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14062_ rbzero.wall_tracer.trackDistY\[-8\] _06786_ _06793_ vssd1 vssd1 vccd1 vccd1
+ _00431_ sky130_fd_sc_hd__o21a_1
XFILLER_113_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11274_ _04051_ _04058_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__nor2_1
XFILLER_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13013_ _05747_ _05769_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__nand2_1
X_10225_ rbzero.tex_g0\[22\] rbzero.tex_g0\[21\] _03166_ vssd1 vssd1 vccd1 vccd1 _03173_
+ sky130_fd_sc_hd__mux2_1
XFILLER_106_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18870_ _04020_ _03464_ _04046_ _02699_ _02334_ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__o41a_1
X_19133__297 clknet_1_0__leaf__02745_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__inv_2
X_17821_ _02073_ _02074_ _02084_ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__a21o_1
XFILLER_79_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10156_ _03136_ vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17752_ _01996_ _02005_ _01992_ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__o21a_1
X_10087_ _03100_ vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__clkbuf_1
X_14964_ _07651_ _07624_ vssd1 vssd1 vccd1 vccd1 _07652_ sky130_fd_sc_hd__nor2_1
X_16703_ _09309_ _09310_ _09311_ vssd1 vssd1 vccd1 vccd1 _09312_ sky130_fd_sc_hd__or3_1
X_13915_ _06661_ _06662_ _06663_ _05265_ _06668_ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__a221o_2
XFILLER_130_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17683_ _01955_ _01956_ _03486_ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__a21oi_1
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14895_ _07549_ _07580_ _07582_ vssd1 vssd1 vccd1 vccd1 _07583_ sky130_fd_sc_hd__nor3_1
X_19422_ rbzero.debug_overlay.vplaneX\[-9\] rbzero.wall_tracer.rayAddendX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__or2_1
X_16634_ _09226_ _09242_ vssd1 vssd1 vccd1 vccd1 _09243_ sky130_fd_sc_hd__xnor2_1
X_13846_ _05367_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__buf_2
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19353_ rbzero.traced_texa\[4\] rbzero.texV\[4\] vssd1 vssd1 vccd1 vccd1 _02835_
+ sky130_fd_sc_hd__nand2_1
X_16565_ _09153_ _09174_ vssd1 vssd1 vccd1 vccd1 _09175_ sky130_fd_sc_hd__xnor2_2
XFILLER_16_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13777_ _05805_ _06071_ _06520_ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__o21bai_1
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10989_ rbzero.row_render.size\[6\] _03774_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__and2_1
XFILLER_90_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18384__28 clknet_1_1__leaf__02434_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__inv_2
X_18304_ _02385_ vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__clkbuf_1
X_15516_ _08072_ _08198_ vssd1 vssd1 vccd1 vccd1 _08200_ sky130_fd_sc_hd__or2_1
XFILLER_149_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12728_ _05467_ _05483_ _05484_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__a21oi_2
X_19284_ rbzero.traced_texa\[-7\] rbzero.texV\[-7\] vssd1 vssd1 vccd1 vccd1 _02777_
+ sky130_fd_sc_hd__nor2_1
X_16496_ _07865_ _08333_ _08978_ _08976_ vssd1 vssd1 vccd1 vccd1 _09106_ sky130_fd_sc_hd__o31a_1
XFILLER_31_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18235_ _02334_ _02344_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__and2_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15447_ _07617_ _07646_ _07756_ _07757_ vssd1 vssd1 vccd1 vccd1 _08132_ sky130_fd_sc_hd__or4_1
X_12659_ _05408_ _05413_ _05415_ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__a21bo_1
XFILLER_175_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18166_ _04828_ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__clkbuf_4
XFILLER_117_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15378_ _08061_ _08051_ _08062_ vssd1 vssd1 vccd1 vccd1 _08063_ sky130_fd_sc_hd__o21ai_2
X_17117_ _09633_ _09654_ vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__or2b_1
XFILLER_129_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14329_ _07016_ _06980_ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18097_ _02253_ vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17048_ _09651_ _09652_ vssd1 vssd1 vccd1 vccd1 _09653_ sky130_fd_sc_hd__nor2_1
XFILLER_172_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__02737_ _02737_ vssd1 vssd1 vccd1 vccd1 clknet_0__02737_ sky130_fd_sc_hd__clkbuf_16
X_09870_ _02986_ vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__clkbuf_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20326_ net386 _01257_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20257_ net317 _01188_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10010_ _03059_ vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09999_ rbzero.tex_r0\[1\] rbzero.tex_r0\[0\] _03050_ vssd1 vssd1 vccd1 vccd1 _03054_
+ sky130_fd_sc_hd__mux2_1
X_20188_ net248 _01119_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[35\] sky130_fd_sc_hd__dfxtp_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ _03474_ _04730_ _04734_ net29 vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__a211oi_1
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10912_ rbzero.tex_r0\[19\] _03696_ _03697_ vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__and3_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ _06410_ _06453_ _06454_ _06456_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__a22o_1
XFILLER_17_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14680_ _07365_ _07367_ _07363_ vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__a21oi_1
X_11892_ _03782_ _04665_ _04666_ _03865_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__a22o_1
Xclkbuf_1_0__f__02726_ clknet_0__02726_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02726_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13631_ _06385_ _06386_ _06387_ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__and3_1
X_10843_ rbzero.row_render.texu\[4\] rbzero.row_render.texu\[3\] _03627_ _03628_ vssd1
+ vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__or4_1
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13562_ _06313_ _06314_ _06317_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__nand3_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16350_ _08836_ _08839_ vssd1 vssd1 vccd1 vccd1 _08962_ sky130_fd_sc_hd__nand2_1
X_10774_ rbzero.traced_texVinit\[5\] rbzero.spi_registers.vshift\[2\] vssd1 vssd1
+ vccd1 vccd1 _03560_ sky130_fd_sc_hd__nor2_1
XFILLER_9_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15301_ _07978_ _07986_ vssd1 vssd1 vccd1 vccd1 _07987_ sky130_fd_sc_hd__nand2_1
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12513_ _05269_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__clkbuf_4
X_16281_ _08229_ _08130_ _08133_ _07494_ vssd1 vssd1 vccd1 vccd1 _08893_ sky130_fd_sc_hd__o22a_1
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13493_ _06241_ _06243_ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__nand2_1
XFILLER_185_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18020_ rbzero.pov.spi_buffer\[62\] rbzero.pov.ready_buffer\[62\] _02208_ vssd1 vssd1
+ vccd1 vccd1 _02212_ sky130_fd_sc_hd__mux2_1
XFILLER_157_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15232_ _07850_ _07918_ vssd1 vssd1 vccd1 vccd1 _07919_ sky130_fd_sc_hd__xnor2_1
X_12444_ _05146_ _05200_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__xor2_2
XFILLER_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15163_ _07793_ _07849_ vssd1 vssd1 vccd1 vccd1 _07850_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12375_ _05097_ _05099_ _05105_ _05127_ _05131_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__a2111o_1
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14114_ _06821_ vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__clkbuf_1
X_11326_ rbzero.debug_overlay.vplaneY\[-7\] _04083_ _04110_ vssd1 vssd1 vccd1 vccd1
+ _04111_ sky130_fd_sc_hd__a21o_1
XFILLER_181_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19971_ net200 _00902_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[51\] sky130_fd_sc_hd__dfxtp_1
X_15094_ _07331_ _07334_ vssd1 vssd1 vccd1 vccd1 _07782_ sky130_fd_sc_hd__and2_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14045_ _06774_ _05373_ _06745_ vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__and3_1
X_19215__372 clknet_1_1__leaf__02752_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__inv_2
X_11257_ _03511_ _03473_ _03781_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__and3b_1
XFILLER_141_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10208_ rbzero.tex_g0\[30\] rbzero.tex_g0\[29\] _03155_ vssd1 vssd1 vccd1 vccd1 _03164_
+ sky130_fd_sc_hd__mux2_1
X_18853_ rbzero.debug_overlay.vplaneY\[-1\] _02637_ vssd1 vssd1 vccd1 vccd1 _02689_
+ sky130_fd_sc_hd__or2_1
XFILLER_67_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11188_ rbzero.tex_r1\[11\] _03664_ _03972_ _03677_ vssd1 vssd1 vccd1 vccd1 _03973_
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17804_ _02056_ _02057_ _02059_ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__and3_1
X_10139_ _03127_ vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__clkbuf_1
X_18784_ rbzero.debug_overlay.facingX\[0\] _02638_ vssd1 vssd1 vccd1 vccd1 _02652_
+ sky130_fd_sc_hd__or2_1
X_15996_ _08325_ _08608_ _08609_ vssd1 vssd1 vccd1 vccd1 _08610_ sky130_fd_sc_hd__o21a_1
XFILLER_48_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17735_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.debug_overlay.vplaneX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__xor2_1
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14947_ _07615_ _07629_ _07634_ vssd1 vssd1 vccd1 vccd1 _07635_ sky130_fd_sc_hd__o21a_1
XFILLER_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17666_ rbzero.wall_tracer.rayAddendX\[-4\] _08463_ _01938_ _01941_ vssd1 vssd1 vccd1
+ vccd1 _00627_ sky130_fd_sc_hd__a22o_1
X_14878_ _07564_ _07565_ vssd1 vssd1 vccd1 vccd1 _07566_ sky130_fd_sc_hd__nor2_1
XFILLER_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19405_ gpout0.clk_div\[0\] net61 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__nor2_1
X_16617_ _09224_ _09225_ vssd1 vssd1 vccd1 vccd1 _09226_ sky130_fd_sc_hd__or2_1
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13829_ _06584_ _06585_ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__nor2_1
XFILLER_23_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17597_ _01880_ _01881_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__nand2_1
XFILLER_51_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19336_ _02816_ _02817_ _02818_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__a21o_1
X_16548_ _09156_ _09157_ vssd1 vssd1 vccd1 vccd1 _09158_ sky130_fd_sc_hd__nor2_1
XFILLER_189_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19267_ rbzero.traced_texa\[-10\] rbzero.texV\[-10\] vssd1 vssd1 vccd1 vccd1 _02763_
+ sky130_fd_sc_hd__or2_1
X_16479_ _08967_ _09075_ vssd1 vssd1 vccd1 vccd1 _09089_ sky130_fd_sc_hd__or2b_1
XFILLER_149_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18218_ _02323_ _02332_ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__and2_1
XFILLER_176_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19198_ clknet_1_0__leaf__02743_ vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__buf_1
XFILLER_15_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18149_ rbzero.spi_registers.got_new_mapd _02261_ vssd1 vssd1 vccd1 vccd1 _02291_
+ sky130_fd_sc_hd__and2_1
XFILLER_191_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20111_ clknet_leaf_90_i_clk _01042_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_116_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09922_ _03013_ vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09853_ _02975_ vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20042_ clknet_leaf_6_i_clk _00973_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09784_ _02939_ vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10490_ _03311_ vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12160_ _04881_ _04921_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__nand2_1
XFILLER_162_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11111_ _03888_ _03889_ _03892_ _03895_ _03896_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__a41o_1
XFILLER_190_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20309_ net369 _01240_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_122_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12091_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__nor2_1
XFILLER_150_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11042_ rbzero.floor_leak\[5\] _03718_ _03685_ rbzero.floor_leak\[4\] _03827_ vssd1
+ vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__o221a_1
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15850_ _03369_ _07825_ _08479_ vssd1 vssd1 vccd1 vccd1 _08480_ sky130_fd_sc_hd__o21a_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ _06865_ _06993_ vssd1 vssd1 vccd1 vccd1 _07489_ sky130_fd_sc_hd__nor2_1
XFILLER_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _08452_ vssd1 vssd1 vccd1 vccd1 _08453_ sky130_fd_sc_hd__buf_4
XFILLER_91_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12993_ _05746_ _05748_ _05749_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__a21o_1
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ _01803_ _01804_ _01810_ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__a21o_1
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14732_ _07416_ _07404_ _07418_ vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__and3_1
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11944_ _04682_ _04712_ _04715_ _04718_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__a211o_1
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__or2_1
X_11875_ _04647_ _04650_ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__nor2_1
XFILLER_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14663_ _06933_ _06939_ vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__nor2_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16402_ _09011_ _09012_ vssd1 vssd1 vccd1 vccd1 _09013_ sky130_fd_sc_hd__xnor2_1
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10826_ _03611_ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__buf_6
X_13614_ _06367_ _06370_ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__or2b_1
X_17382_ _01685_ vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__clkbuf_1
X_14594_ _07007_ _07281_ _07249_ _07248_ vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__o31a_1
XFILLER_38_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19121_ clknet_1_1__leaf__02743_ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__buf_1
X_16333_ _08763_ _08820_ _08944_ vssd1 vssd1 vccd1 vccd1 _08945_ sky130_fd_sc_hd__a21oi_1
X_10757_ rbzero.traced_texVinit\[4\] rbzero.spi_registers.vshift\[1\] vssd1 vssd1
+ vccd1 vccd1 _03543_ sky130_fd_sc_hd__or2_1
X_13545_ _06295_ _06301_ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__or2_1
XFILLER_158_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16264_ _08749_ _08752_ _08874_ vssd1 vssd1 vccd1 vccd1 _08876_ sky130_fd_sc_hd__and3_1
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13476_ _06072_ _06157_ vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__or2_1
XFILLER_145_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10688_ _03479_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__buf_2
XFILLER_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18003_ rbzero.pov.spi_buffer\[54\] rbzero.pov.ready_buffer\[54\] _02197_ vssd1 vssd1
+ vccd1 vccd1 _02203_ sky130_fd_sc_hd__mux2_1
X_15215_ _07899_ _07901_ vssd1 vssd1 vccd1 vccd1 _07902_ sky130_fd_sc_hd__and2b_1
X_12427_ _05161_ _05183_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__xor2_1
X_16195_ _08802_ _08807_ vssd1 vssd1 vccd1 vccd1 _08808_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15146_ _07726_ _07704_ vssd1 vssd1 vccd1 vccd1 _07833_ sky130_fd_sc_hd__or2b_1
X_12358_ rbzero.wall_tracer.visualWallDist\[-11\] rbzero.wall_tracer.rayAddendY\[-3\]
+ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__mux2_1
XFILLER_126_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11309_ rbzero.debug_overlay.facingY\[-3\] _04092_ _04093_ rbzero.debug_overlay.facingY\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__a22o_1
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19954_ net183 _00885_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[34\] sky130_fd_sc_hd__dfxtp_1
X_15077_ _07761_ vssd1 vssd1 vccd1 vccd1 _07765_ sky130_fd_sc_hd__inv_2
X_12289_ _05038_ _05039_ _05044_ _05045_ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__o31ai_4
X_14028_ rbzero.wall_tracer.stepDistY\[6\] _06767_ _06718_ vssd1 vssd1 vccd1 vccd1
+ _06768_ sky130_fd_sc_hd__mux2_1
XFILLER_171_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19885_ clknet_leaf_21_i_clk _00816_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18836_ rbzero.pov.ready_buffer\[21\] _02663_ _02680_ _02672_ vssd1 vssd1 vccd1 vccd1
+ _01058_ sky130_fd_sc_hd__o211a_1
XFILLER_45_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__02436_ _02436_ vssd1 vssd1 vccd1 vccd1 clknet_0__02436_ sky130_fd_sc_hd__clkbuf_16
X_18767_ rbzero.pov.ready_buffer\[35\] _02636_ _02641_ _02586_ vssd1 vssd1 vccd1 vccd1
+ _01028_ sky130_fd_sc_hd__o211a_1
XFILLER_55_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15979_ rbzero.wall_tracer.trackDistX\[0\] rbzero.wall_tracer.stepDistX\[0\] vssd1
+ vssd1 vccd1 vccd1 _08593_ sky130_fd_sc_hd__nor2_1
X_17718_ _01986_ _01987_ _01988_ _01974_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__a211o_1
X_18698_ rbzero.pov.ready_buffer\[45\] vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__inv_2
X_17649_ rbzero.debug_overlay.vplaneX\[-7\] rbzero.wall_tracer.rayAddendX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__nand2_1
XFILLER_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19319_ rbzero.traced_texa\[-1\] rbzero.texV\[-1\] vssd1 vssd1 vccd1 vccd1 _02806_
+ sky130_fd_sc_hd__and2_1
XFILLER_149_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09905_ _03004_ vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20025_ clknet_leaf_87_i_clk _00956_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09836_ rbzero.tex_r1\[12\] rbzero.tex_r1\[13\] _02965_ vssd1 vssd1 vccd1 vccd1 _02967_
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09767_ _02930_ vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11660_ _03689_ _04436_ _04440_ _03679_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__a211o_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _03353_ _03369_ rbzero.map_rom.i_col\[4\] _03406_ vssd1 vssd1 vccd1 vccd1
+ _03407_ sky130_fd_sc_hd__or4_1
XFILLER_179_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11591_ _04370_ _04371_ _04372_ _04192_ _04179_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__o221a_1
X_13330_ _06060_ _06086_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__xnor2_2
XFILLER_195_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10542_ _03338_ vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__buf_6
XFILLER_109_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13261_ _05964_ _06014_ _06016_ _06017_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__or4_1
X_10473_ rbzero.tex_b0\[32\] rbzero.tex_b0\[31\] _03302_ vssd1 vssd1 vccd1 vccd1 _03303_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15000_ _07645_ _07686_ _07687_ vssd1 vssd1 vccd1 vccd1 _07688_ sky130_fd_sc_hd__o21ai_1
X_12212_ rbzero.wall_tracer.trackDistY\[-8\] vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__inv_2
XFILLER_108_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13192_ _05907_ _05948_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__xor2_1
XFILLER_109_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12143_ _04899_ _04866_ _04853_ _04848_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__a211o_1
XFILLER_150_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16951_ _09555_ _09556_ vssd1 vssd1 vccd1 vccd1 _09557_ sky130_fd_sc_hd__and2b_1
X_12074_ rbzero.wall_tracer.state\[6\] vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__inv_4
XFILLER_96_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11025_ rbzero.row_render.size\[1\] _03809_ _03810_ _03771_ vssd1 vssd1 vccd1 vccd1
+ _03811_ sky130_fd_sc_hd__a31o_1
X_15902_ _08524_ _07817_ vssd1 vssd1 vccd1 vccd1 _08525_ sky130_fd_sc_hd__and2_1
X_19670_ clknet_leaf_11_i_clk _00601_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f1 sky130_fd_sc_hd__dfxtp_1
XFILLER_103_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16882_ _09021_ _09035_ vssd1 vssd1 vccd1 vccd1 _09489_ sky130_fd_sc_hd__nor2_1
X_18621_ rbzero.pov.sclk_buffer\[1\] rbzero.pov.sclk_buffer\[0\] _04827_ vssd1 vssd1
+ vccd1 vccd1 _02530_ sky130_fd_sc_hd__mux2_1
XFILLER_77_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15833_ rbzero.wall_tracer.wall\[0\] rbzero.row_render.wall\[0\] _08464_ vssd1 vssd1
+ vccd1 vccd1 _08465_ sky130_fd_sc_hd__mux2_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18552_ _02494_ vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _04040_ _08438_ vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__nor2_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _05709_ _05710_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__xor2_1
XFILLER_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19026__201 clknet_1_1__leaf__02734_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__inv_2
XFILLER_166_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ _01777_ _01794_ vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__xnor2_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14715_ _07400_ _07402_ vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__xnor2_1
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18483_ _02458_ vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11927_ _04672_ net62 vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__or2_1
X_15695_ _07992_ _08252_ _08251_ vssd1 vssd1 vccd1 vccd1 _08378_ sky130_fd_sc_hd__or3_1
XFILLER_60_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17434_ _01726_ _01727_ _01729_ _01730_ _03497_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__o311a_1
X_14646_ _07011_ _07333_ vssd1 vssd1 vccd1 vccd1 _07334_ sky130_fd_sc_hd__nor2_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11858_ net47 _04626_ _04627_ _04633_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__a22o_1
XFILLER_33_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10809_ _03593_ _03594_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__nor2_1
XANTENNA_19 rbzero.debug_overlay.facingX\[-1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17365_ rbzero.spi_registers.new_mapd\[11\] rbzero.spi_registers.spi_buffer\[11\]
+ _01662_ vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__mux2_1
XFILLER_186_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14577_ _07049_ vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__clkbuf_4
XFILLER_14_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11789_ net16 net15 vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__nor2_1
XFILLER_13_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16316_ _08802_ _08807_ _08805_ vssd1 vssd1 vccd1 vccd1 _08928_ sky130_fd_sc_hd__a21boi_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13528_ _06278_ _06280_ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__or2_1
XFILLER_9_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17296_ rbzero.wall_tracer.trackDistY\[5\] rbzero.wall_tracer.stepDistY\[5\] vssd1
+ vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__and2_1
XFILLER_12_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16247_ _07856_ _08316_ vssd1 vssd1 vccd1 vccd1 _08859_ sky130_fd_sc_hd__and2_1
X_13459_ _06212_ _06214_ vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__nand2_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16178_ _08789_ _08790_ vssd1 vssd1 vccd1 vccd1 _08791_ sky130_fd_sc_hd__nor2_1
XFILLER_103_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19072__243 clknet_1_0__leaf__02738_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__inv_2
XFILLER_141_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15129_ _07696_ _07698_ vssd1 vssd1 vccd1 vccd1 _07817_ sky130_fd_sc_hd__xor2_4
XFILLER_114_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_92_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_114_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19937_ net166 _00868_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__04486_ clknet_0__04486_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04486_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_130_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19868_ clknet_leaf_24_i_clk _00799_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18819_ rbzero.debug_overlay.vplaneX\[-6\] _02660_ vssd1 vssd1 vccd1 vccd1 _02671_
+ sky130_fd_sc_hd__or2_1
XFILLER_56_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19799_ clknet_leaf_16_i_clk _00730_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_83_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_30_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_45_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20008_ clknet_leaf_75_i_clk _00939_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09819_ rbzero.tex_r1\[20\] rbzero.tex_r1\[21\] _02954_ vssd1 vssd1 vccd1 vccd1 _02958_
+ sky130_fd_sc_hd__mux2_1
XFILLER_100_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12830_ _05477_ _05480_ _05485_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__and3_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _05516_ _05517_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__or2_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _07181_ _07187_ vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _04487_ _04314_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__nand2_1
XFILLER_188_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15480_ _08162_ _08164_ vssd1 vssd1 vccd1 vccd1 _08165_ sky130_fd_sc_hd__xor2_2
X_12692_ _05210_ _05445_ _05446_ _05323_ _05448_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__a32oi_4
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11643_ rbzero.tex_b1\[49\] rbzero.tex_b1\[48\] _04376_ vssd1 vssd1 vccd1 vccd1 _04424_
+ sky130_fd_sc_hd__mux2_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14431_ _06893_ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__buf_2
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17150_ _01481_ _01493_ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11574_ _04353_ _04354_ _04355_ _04192_ _04179_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__o221a_1
X_14362_ _06985_ _04922_ _07026_ vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__or3_1
Xinput17 i_gpout2_sel[2] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_6
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput28 i_gpout4_sel[1] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_4
X_16101_ _08299_ _08302_ _08430_ _08714_ _08429_ vssd1 vssd1 vccd1 vccd1 _08715_ sky130_fd_sc_hd__a32oi_4
Xinput39 i_mode[0] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_16
XFILLER_168_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10525_ rbzero.tex_b0\[7\] rbzero.tex_b0\[6\] _03324_ vssd1 vssd1 vccd1 vccd1 _03330_
+ sky130_fd_sc_hd__mux2_1
X_13313_ _05905_ _06069_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__or2_1
X_17081_ _09672_ _09685_ vssd1 vssd1 vccd1 vccd1 _09686_ sky130_fd_sc_hd__xor2_1
XFILLER_122_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14293_ rbzero.debug_overlay.playerY\[-3\] _06956_ vssd1 vssd1 vccd1 vccd1 _06981_
+ sky130_fd_sc_hd__nand2_1
XFILLER_196_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16032_ _08229_ _07137_ vssd1 vssd1 vccd1 vccd1 _08646_ sky130_fd_sc_hd__or2_1
XFILLER_157_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13244_ _05593_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__clkbuf_4
X_10456_ rbzero.tex_b0\[40\] rbzero.tex_b0\[39\] _03291_ vssd1 vssd1 vccd1 vccd1 _03294_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ _05927_ _05931_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__and2_1
X_10387_ rbzero.tex_b1\[8\] rbzero.tex_b1\[9\] _03254_ vssd1 vssd1 vccd1 vccd1 _03258_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12126_ _04873_ _04887_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__nor2_1
XFILLER_2_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17983_ _02192_ vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19722_ clknet_leaf_87_i_clk _00653_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16934_ _09007_ _09039_ vssd1 vssd1 vccd1 vccd1 _09540_ sky130_fd_sc_hd__nor2_1
X_12057_ _04827_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__buf_6
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11008_ rbzero.row_render.size\[9\] _03778_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__nand2_1
X_19653_ clknet_leaf_18_i_clk _00584_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16865_ _09283_ _09471_ vssd1 vssd1 vccd1 vccd1 _09472_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18604_ _02521_ vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15816_ rbzero.traced_texa\[-3\] _08461_ _08459_ rbzero.wall_tracer.visualWallDist\[-3\]
+ vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__a22o_1
X_19584_ clknet_leaf_61_i_clk _00515_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16796_ _09208_ _09402_ vssd1 vssd1 vccd1 vccd1 _09404_ sky130_fd_sc_hd__or2_1
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18535_ _02485_ vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__clkbuf_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15747_ _08294_ _08429_ vssd1 vssd1 vccd1 vccd1 _08430_ sky130_fd_sc_hd__xnor2_4
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12959_ _05713_ _05714_ _05715_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__a21oi_1
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18466_ _02449_ vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__clkbuf_1
X_15678_ _08233_ _08359_ _08360_ vssd1 vssd1 vccd1 vccd1 _08361_ sky130_fd_sc_hd__o21ba_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17417_ _08453_ _01713_ _01715_ vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__a21o_1
XFILLER_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14629_ _07308_ _07315_ _07316_ vssd1 vssd1 vccd1 vccd1 _07317_ sky130_fd_sc_hd__a21oi_1
XFILLER_53_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17348_ _01666_ vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17279_ rbzero.wall_tracer.trackDistY\[2\] _01558_ _01608_ _08959_ vssd1 vssd1 vccd1
+ vccd1 _00573_ sky130_fd_sc_hd__o22a_1
XFILLER_162_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20290_ net350 _01221_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18937__121 clknet_1_1__leaf__02725_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__inv_2
XFILLER_161_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18983__163 clknet_1_0__leaf__02729_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__inv_2
XFILLER_169_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19079__249 clknet_1_1__leaf__02739_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__inv_2
XFILLER_193_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10310_ _03217_ vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11290_ _04044_ _04047_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__nand2_1
X_20488_ clknet_leaf_41_i_clk _01419_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10241_ _03181_ vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10172_ _03145_ vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_121_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14980_ _07654_ _07658_ vssd1 vssd1 vccd1 vccd1 _07668_ sky130_fd_sc_hd__xor2_1
XFILLER_87_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13931_ _06601_ _06614_ _06638_ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__o21ai_1
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16650_ _09140_ _09143_ _09139_ vssd1 vssd1 vccd1 vccd1 _09259_ sky130_fd_sc_hd__a21bo_1
XFILLER_75_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13862_ _06615_ _06618_ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__nor2_1
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15601_ _08243_ _08283_ vssd1 vssd1 vccd1 vccd1 _08285_ sky130_fd_sc_hd__or2_1
X_12813_ _05567_ _05568_ _05569_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__o21a_1
XFILLER_16_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16581_ _09189_ _09190_ vssd1 vssd1 vccd1 vccd1 _09191_ sky130_fd_sc_hd__nand2_1
X_13793_ _06383_ _06536_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__or2_1
XFILLER_76_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18320_ _02394_ vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__clkbuf_1
X_15532_ _08214_ _08215_ vssd1 vssd1 vccd1 vccd1 _08216_ sky130_fd_sc_hd__nor2_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _05487_ _05500_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__and2b_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18251_ rbzero.spi_registers.new_vshift\[4\] _02348_ _02354_ _02314_ vssd1 vssd1
+ vccd1 vccd1 _00799_ sky130_fd_sc_hd__o211a_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _08143_ _08146_ _08138_ vssd1 vssd1 vccd1 vccd1 _08148_ sky130_fd_sc_hd__a21oi_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _05316_ _05332_ _05375_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__mux2_1
X_17202_ rbzero.wall_tracer.trackDistY\[-8\] rbzero.wall_tracer.stepDistY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__nand2_1
XFILLER_187_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14414_ rbzero.wall_tracer.stepDistX\[0\] vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__inv_2
X_11626_ rbzero.tex_b1\[39\] rbzero.tex_b1\[38\] _03617_ vssd1 vssd1 vccd1 vccd1 _04407_
+ sky130_fd_sc_hd__mux2_1
X_18182_ rbzero.mapdyw\[1\] _02291_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__or2_1
X_15394_ _06979_ _07007_ _07332_ _07786_ vssd1 vssd1 vccd1 vccd1 _08079_ sky130_fd_sc_hd__or4_1
XFILLER_156_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17133_ _09658_ _09689_ _09687_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__a21bo_1
X_19138__302 clknet_1_1__leaf__02745_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__inv_2
XFILLER_11_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14345_ rbzero.debug_overlay.playerX\[-2\] _06987_ rbzero.debug_overlay.playerX\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__o21ai_1
X_11557_ _04336_ _04337_ _04338_ _04192_ _04179_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__o221a_1
XFILLER_129_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17064_ _09666_ _09667_ vssd1 vssd1 vccd1 vccd1 _09669_ sky130_fd_sc_hd__and2_1
XFILLER_156_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10508_ rbzero.tex_b0\[15\] rbzero.tex_b0\[14\] _03313_ vssd1 vssd1 vccd1 vccd1 _03321_
+ sky130_fd_sc_hd__mux2_1
X_11488_ _04268_ _04269_ _04270_ _03917_ _03674_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__o221a_1
X_14276_ _06887_ _06963_ vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__or2_1
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16015_ _08627_ _08628_ vssd1 vssd1 vccd1 vccd1 _08629_ sky130_fd_sc_hd__nor2_1
X_10439_ rbzero.tex_b0\[48\] rbzero.tex_b0\[47\] _03280_ vssd1 vssd1 vccd1 vccd1 _03285_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__02753_ _02753_ vssd1 vssd1 vccd1 vccd1 clknet_0__02753_ sky130_fd_sc_hd__clkbuf_16
X_13227_ _05982_ _05983_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__nor2_2
XFILLER_100_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13158_ _05609_ _05593_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__nor2_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ rbzero.debug_overlay.facingY\[-1\] rbzero.wall_tracer.rayAddendY\[7\] vssd1
+ vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__nor2_1
X_13089_ _05834_ _05845_ _05832_ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__and3b_1
X_17966_ _02183_ vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19705_ clknet_leaf_71_i_clk _00636_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_16917_ _09417_ _09419_ _09418_ vssd1 vssd1 vccd1 vccd1 _09524_ sky130_fd_sc_hd__o21ba_1
X_17897_ _02147_ vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19184__344 clknet_1_0__leaf__02749_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__inv_2
XFILLER_66_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16848_ _09335_ _09344_ _09342_ vssd1 vssd1 vccd1 vccd1 _09455_ sky130_fd_sc_hd__a21oi_1
XFILLER_38_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19636_ clknet_leaf_60_i_clk _00567_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19567_ clknet_leaf_36_i_clk _00498_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_81_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16779_ _09279_ _09283_ _09280_ vssd1 vssd1 vccd1 vccd1 _09387_ sky130_fd_sc_hd__a21boi_1
XFILLER_80_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18518_ _02476_ vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__clkbuf_1
X_19498_ clknet_leaf_46_i_clk _00444_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[5\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18449_ clknet_1_0__leaf__02440_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__buf_1
XFILLER_178_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20411_ net471 _01342_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20342_ net402 _01273_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20273_ net333 _01204_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__02742_ clknet_0__02742_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02742_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10790_ _03572_ _03575_ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__nor2_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12460_ _05105_ _05216_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__xnor2_4
XFILLER_138_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11411_ rbzero.tex_g0\[50\] _03727_ _03652_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__a21o_1
XFILLER_166_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_73 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_73/HI o_rgb[0] sky130_fd_sc_hd__conb_1
XFILLER_32_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12391_ rbzero.wall_tracer.visualWallDist\[3\] _03479_ vssd1 vssd1 vccd1 vccd1 _05148_
+ sky130_fd_sc_hd__nor2_1
Xtop_ew_algofoogle_84 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_84/HI o_rgb[13] sky130_fd_sc_hd__conb_1
XFILLER_32_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_95 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_95/HI zeros[4] sky130_fd_sc_hd__conb_1
XFILLER_125_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11342_ rbzero.debug_overlay.playerX\[-7\] _04083_ _04085_ rbzero.debug_overlay.playerX\[-5\]
+ _04126_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__a221o_1
X_14130_ rbzero.wall_tracer.stepDistX\[2\] _06746_ _06825_ vssd1 vssd1 vccd1 vccd1
+ _06830_ sky130_fd_sc_hd__mux2_1
XFILLER_126_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11273_ _03460_ _04057_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__or2_1
X_14061_ rbzero.wall_tracer.visualWallDist\[-8\] _03496_ _06791_ rbzero.wall_tracer.trackDistX\[-8\]
+ _03485_ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__o221a_1
XFILLER_165_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10224_ _03172_ vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__clkbuf_1
X_13012_ _05516_ _05503_ _05768_ _05697_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17820_ _02081_ _02070_ _02083_ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__a21oi_1
XFILLER_95_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10155_ rbzero.tex_g0\[55\] rbzero.tex_g0\[54\] _03132_ vssd1 vssd1 vccd1 vccd1 _03136_
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17751_ _02018_ _02019_ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__and2b_1
XFILLER_43_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10086_ rbzero.tex_g1\[23\] rbzero.tex_g1\[24\] _03095_ vssd1 vssd1 vccd1 vccd1 _03100_
+ sky130_fd_sc_hd__mux2_1
X_14963_ _07625_ vssd1 vssd1 vccd1 vccd1 _07651_ sky130_fd_sc_hd__inv_2
XFILLER_48_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16702_ _09199_ _09201_ _09198_ vssd1 vssd1 vccd1 vccd1 _09311_ sky130_fd_sc_hd__a21boi_1
X_13914_ _05476_ _06667_ _06630_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__a21o_1
X_17682_ _01951_ _01952_ _01954_ vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__o21ai_1
X_14894_ _06873_ _07581_ _07530_ _06866_ vssd1 vssd1 vccd1 vccd1 _07582_ sky130_fd_sc_hd__o22a_1
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19421_ _02878_ _02879_ rbzero.wall_tracer.rayAddendY\[-6\] _08449_ vssd1 vssd1 vccd1
+ vccd1 _01444_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16633_ _09240_ _09241_ vssd1 vssd1 vccd1 vccd1 _09242_ sky130_fd_sc_hd__xor2_1
X_13845_ _06598_ _06600_ _06601_ vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__mux2_1
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19352_ rbzero.traced_texa\[4\] rbzero.texV\[4\] vssd1 vssd1 vccd1 vccd1 _02834_
+ sky130_fd_sc_hd__or2_1
XFILLER_188_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16564_ _09172_ _09173_ vssd1 vssd1 vccd1 vccd1 _09174_ sky130_fd_sc_hd__xor2_2
X_13776_ _05805_ _06156_ _06532_ vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__or3_1
XFILLER_200_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10988_ rbzero.row_render.size\[5\] rbzero.row_render.size\[4\] _03773_ vssd1 vssd1
+ vccd1 vccd1 _03774_ sky130_fd_sc_hd__or3_1
X_18303_ rbzero.spi_registers.spi_buffer\[5\] rbzero.spi_registers.new_leak\[5\] _02379_
+ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__mux2_1
X_15515_ _08072_ _08198_ vssd1 vssd1 vccd1 vccd1 _08199_ sky130_fd_sc_hd__nand2_1
XFILLER_128_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12727_ _05449_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__clkbuf_4
X_19283_ rbzero.texV\[-8\] _02675_ _02709_ _02776_ vssd1 vssd1 vccd1 vccd1 _01409_
+ sky130_fd_sc_hd__a22o_1
X_16495_ _09100_ _09104_ vssd1 vssd1 vccd1 vccd1 _09105_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18234_ rbzero.color_floor\[4\] rbzero.spi_registers.new_floor\[4\] _02335_ vssd1
+ vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__mux2_1
XFILLER_31_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15446_ _07877_ _08130_ vssd1 vssd1 vccd1 vccd1 _08131_ sky130_fd_sc_hd__nor2_1
X_12658_ _05414_ _05339_ _05342_ _05209_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__o31a_1
XFILLER_169_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18165_ rbzero.map_overlay.i_mapdy\[1\] _02292_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__or2_1
X_11609_ _03896_ _04390_ _03518_ _03529_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__or4bb_1
XFILLER_156_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15377_ _07940_ _08047_ vssd1 vssd1 vccd1 vccd1 _08062_ sky130_fd_sc_hd__nand2_1
XFILLER_50_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12589_ _05344_ _05345_ _05338_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__mux2_1
XFILLER_117_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17116_ _09691_ _09692_ _01459_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__o21a_1
XFILLER_190_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14328_ rbzero.debug_overlay.playerY\[-2\] vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__inv_2
XFILLER_117_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18096_ rbzero.spi_registers.ss_buffer\[1\] rbzero.spi_registers.ss_buffer\[0\] _04834_
+ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__mux2_1
XFILLER_183_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17047_ _09635_ _09650_ vssd1 vssd1 vccd1 vccd1 _09652_ sky130_fd_sc_hd__nor2_1
XFILLER_144_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14259_ _06887_ _06946_ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__or2_1
XFILLER_143_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__02736_ _02736_ vssd1 vssd1 vccd1 vccd1 clknet_0__02736_ sky130_fd_sc_hd__clkbuf_16
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18998_ clknet_1_1__leaf__02440_ vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__buf_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17949_ _02174_ vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19619_ clknet_leaf_52_i_clk _00550_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18907__94 clknet_1_0__leaf__02441_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__inv_2
XFILLER_55_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20325_ net385 _01256_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20256_ net316 _01187_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20187_ net247 _01118_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09998_ _03053_ vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_130_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ _03782_ _04731_ _04732_ _03865_ _04733_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__a221o_1
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10911_ _03613_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__buf_4
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02725_ clknet_0__02725_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02725_
+ sky130_fd_sc_hd__clkbuf_16
X_11891_ net22 net21 vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__and2_1
XFILLER_151_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13630_ _06103_ _06071_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__nor2_1
XFILLER_71_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10842_ rbzero.row_render.texu\[2\] rbzero.row_render.texu\[1\] vssd1 vssd1 vccd1
+ vccd1 _03628_ sky130_fd_sc_hd__nand2_1
XFILLER_71_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13561_ _06313_ _06314_ _06317_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__a21o_1
X_10773_ rbzero.traced_texVinit\[5\] rbzero.spi_registers.vshift\[2\] vssd1 vssd1
+ vccd1 vccd1 _03559_ sky130_fd_sc_hd__and2_1
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15300_ _07983_ _07985_ vssd1 vssd1 vccd1 vccd1 _07986_ sky130_fd_sc_hd__xor2_1
XFILLER_9_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12512_ _05268_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__buf_2
XFILLER_197_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16280_ _08229_ _08133_ _08773_ vssd1 vssd1 vccd1 vccd1 _08892_ sky130_fd_sc_hd__or3_1
XFILLER_200_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13492_ _06149_ _06245_ _06246_ _06248_ vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__a22oi_2
XFILLER_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15231_ _07916_ _07917_ vssd1 vssd1 vccd1 vccd1 _07918_ sky130_fd_sc_hd__and2b_1
XFILLER_138_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12443_ _05199_ _05133_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__nand2_2
XFILLER_200_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15162_ _07847_ _07848_ vssd1 vssd1 vccd1 vccd1 _07849_ sky130_fd_sc_hd__nor2_1
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12374_ _03487_ _05128_ _05129_ _05130_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_176_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14113_ rbzero.wall_tracer.stepDistX\[-6\] _06686_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _06821_ sky130_fd_sc_hd__mux2_1
XFILLER_125_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11325_ rbzero.debug_overlay.vplaneY\[-9\] _04081_ _04084_ rbzero.debug_overlay.vplaneY\[-6\]
+ _03854_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__a221o_1
X_19970_ net199 _00901_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15093_ _07289_ _07262_ vssd1 vssd1 vccd1 vccd1 _07781_ sky130_fd_sc_hd__or2b_1
XFILLER_181_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18921_ clknet_1_0__leaf__02440_ vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__buf_1
X_11256_ gpout0.hpos\[4\] _04040_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__nor2_1
X_14044_ _06780_ vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ _03163_ vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11187_ rbzero.tex_r1\[10\] _03620_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__or2_1
X_18852_ rbzero.pov.ready_buffer\[7\] _02666_ _02688_ _02675_ vssd1 vssd1 vccd1 vccd1
+ _01066_ sky130_fd_sc_hd__a211o_1
XFILLER_80_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10138_ rbzero.tex_g0\[63\] rbzero.tex_g0\[62\] _03050_ vssd1 vssd1 vccd1 vccd1 _03127_
+ sky130_fd_sc_hd__mux2_1
X_17803_ _02057_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__inv_2
XFILLER_0_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18783_ rbzero.pov.ready_buffer\[41\] _02644_ _02650_ _02651_ vssd1 vssd1 vccd1 vccd1
+ _01034_ sky130_fd_sc_hd__a211o_1
XFILLER_79_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15995_ _07972_ _07856_ _07959_ _08069_ vssd1 vssd1 vccd1 vccd1 _08609_ sky130_fd_sc_hd__or4_1
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17734_ _01986_ _01990_ _02002_ _02003_ _03486_ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__a311oi_1
X_14946_ _07630_ _07633_ vssd1 vssd1 vccd1 vccd1 _07634_ sky130_fd_sc_hd__nand2_1
X_10069_ rbzero.tex_g1\[31\] rbzero.tex_g1\[32\] _03084_ vssd1 vssd1 vccd1 vccd1 _03091_
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17665_ _01722_ _01939_ _01940_ _08452_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__a31o_1
X_14877_ _07548_ _07563_ vssd1 vssd1 vccd1 vccd1 _07565_ sky130_fd_sc_hd__and2_1
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16616_ _09222_ _09223_ vssd1 vssd1 vccd1 vccd1 _09225_ sky130_fd_sc_hd__and2_1
X_19404_ rbzero.traced_texVinit\[10\] _02868_ _08454_ _08958_ vssd1 vssd1 vccd1 vccd1
+ _01438_ sky130_fd_sc_hd__a22o_1
XFILLER_63_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13828_ _06224_ _06583_ vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__nor2_1
X_17596_ _01786_ rbzero.wall_tracer.rayAddendY\[9\] vssd1 vssd1 vccd1 vccd1 _01881_
+ sky130_fd_sc_hd__nand2_1
XFILLER_51_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16547_ _08245_ _08391_ _08678_ _08247_ vssd1 vssd1 vccd1 vccd1 _09157_ sky130_fd_sc_hd__o22a_1
X_19335_ _02819_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__inv_2
X_13759_ _06337_ _06513_ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__or2_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19266_ _02759_ _02760_ _02761_ _02762_ rbzero.texV\[-11\] vssd1 vssd1 vccd1 vccd1
+ _01406_ sky130_fd_sc_hd__a32o_1
X_16478_ rbzero.wall_tracer.trackDistX\[3\] _08553_ _09081_ _09088_ vssd1 vssd1 vccd1
+ vccd1 _00552_ sky130_fd_sc_hd__o22a_1
X_18217_ rbzero.color_sky\[5\] rbzero.spi_registers.new_sky\[5\] _02320_ vssd1 vssd1
+ vccd1 vccd1 _02332_ sky130_fd_sc_hd__mux2_1
X_15429_ _08096_ _08113_ vssd1 vssd1 vccd1 vccd1 _08114_ sky130_fd_sc_hd__xnor2_1
XFILLER_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18148_ _02289_ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__buf_2
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18079_ _02243_ vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20110_ clknet_leaf_77_i_clk _01041_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
X_09921_ rbzero.tex_r0\[38\] rbzero.tex_r0\[37\] _03006_ vssd1 vssd1 vccd1 vccd1 _03013_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20041_ clknet_leaf_5_i_clk _00972_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_09852_ rbzero.tex_r1\[4\] rbzero.tex_r1\[5\] _02965_ vssd1 vssd1 vccd1 vccd1 _02975_
+ sky130_fd_sc_hd__mux2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ rbzero.tex_r1\[37\] rbzero.tex_r1\[38\] _02932_ vssd1 vssd1 vccd1 vccd1 _02939_
+ sky130_fd_sc_hd__mux2_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__02441_ clknet_0__02441_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02441_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11110_ _03530_ _03532_ _03533_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__or3_2
XFILLER_190_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20308_ net368 _01239_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12090_ _04850_ _04851_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__nor2_1
XFILLER_162_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11041_ rbzero.floor_leak\[3\] _03624_ _03684_ rbzero.floor_leak\[4\] _03826_ vssd1
+ vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__a221o_1
X_20239_ net299 _01170_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_122_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ _07486_ _07481_ vssd1 vssd1 vccd1 vccd1 _07488_ sky130_fd_sc_hd__xor2_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _08451_ vssd1 vssd1 vccd1 vccd1 _08452_ sky130_fd_sc_hd__clkbuf_4
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12992_ _05745_ _05733_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__and2b_1
XFILLER_57_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14731_ _07416_ _07404_ _07418_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__a21oi_1
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ net43 _04668_ _04685_ _04716_ _04717_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__a311o_1
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _08452_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__buf_4
XFILLER_55_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14662_ _07343_ _07349_ vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__xor2_1
X_11874_ _04624_ _04648_ _04649_ _04635_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__a22o_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16401_ _08862_ _07857_ vssd1 vssd1 vccd1 vccd1 _09012_ sky130_fd_sc_hd__nor2_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13613_ _05805_ _06035_ _06367_ _06369_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__or4_1
X_10825_ _03610_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__buf_4
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17381_ _03343_ _01684_ _08507_ vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__mux2_1
X_14593_ _07052_ vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__clkbuf_4
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19120_ clknet_1_1__leaf__04486_ vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__buf_1
X_16332_ _08817_ _08819_ vssd1 vssd1 vccd1 vccd1 _08944_ sky130_fd_sc_hd__nor2_1
XFILLER_198_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13544_ _06247_ _06296_ _06297_ _06300_ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10756_ rbzero.traced_texVinit\[4\] rbzero.spi_registers.vshift\[1\] vssd1 vssd1
+ vccd1 vccd1 _03542_ sky130_fd_sc_hd__nand2_1
XFILLER_41_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16263_ _08749_ _08752_ _08874_ vssd1 vssd1 vccd1 vccd1 _08875_ sky130_fd_sc_hd__a21oi_1
XFILLER_125_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13475_ _05990_ _06156_ _06231_ vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__nor3_2
XFILLER_201_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10687_ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__clkbuf_4
X_18002_ _02202_ vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__clkbuf_1
X_15214_ _07199_ _07757_ _07900_ vssd1 vssd1 vccd1 vccd1 _07901_ sky130_fd_sc_hd__o21bai_1
XFILLER_139_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12426_ _05159_ _05157_ _05153_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__a21oi_2
XFILLER_199_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16194_ _08806_ vssd1 vssd1 vccd1 vccd1 _08807_ sky130_fd_sc_hd__buf_2
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15145_ _07703_ _07807_ _07831_ vssd1 vssd1 vccd1 vccd1 _07832_ sky130_fd_sc_hd__a21oi_2
X_12357_ _05110_ _05111_ _05113_ _05072_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__o22a_2
XFILLER_114_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ _03782_ _04051_ _04057_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__nor3_4
XFILLER_114_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19953_ net182 _00884_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[33\] sky130_fd_sc_hd__dfxtp_1
X_15076_ _07746_ _07763_ vssd1 vssd1 vccd1 vccd1 _07764_ sky130_fd_sc_hd__xnor2_2
XFILLER_142_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12288_ rbzero.debug_overlay.facingX\[-6\] rbzero.wall_tracer.rayAddendX\[2\] vssd1
+ vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__nand2_1
XFILLER_141_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14027_ _05373_ _06715_ _06744_ _06763_ _06630_ vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__a221o_2
X_11239_ gpout0.vpos\[5\] _03523_ _03524_ _03517_ _04023_ vssd1 vssd1 vccd1 vccd1
+ _04024_ sky130_fd_sc_hd__a221o_1
X_19884_ clknet_leaf_18_i_clk _00815_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_floor
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18931__116 clknet_1_1__leaf__02724_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__inv_2
X_18835_ _02094_ _02635_ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__nand2_1
XFILLER_1_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__02435_ _02435_ vssd1 vssd1 vccd1 vccd1 clknet_0__02435_ sky130_fd_sc_hd__clkbuf_16
XFILLER_83_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18766_ rbzero.debug_overlay.facingX\[-7\] _02638_ vssd1 vssd1 vccd1 vccd1 _02641_
+ sky130_fd_sc_hd__or2_1
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15978_ _04966_ _07102_ vssd1 vssd1 vccd1 vccd1 _08592_ sky130_fd_sc_hd__nor2_1
XFILLER_95_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14929_ _07119_ vssd1 vssd1 vccd1 vccd1 _07617_ sky130_fd_sc_hd__buf_2
X_17717_ _01972_ rbzero.wall_tracer.rayAddendX\[0\] _01971_ vssd1 vssd1 vccd1 vccd1
+ _01988_ sky130_fd_sc_hd__o21a_1
XFILLER_36_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18697_ _02587_ vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__buf_2
XFILLER_36_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17648_ _01921_ _01924_ _01922_ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__o21a_1
XFILLER_64_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17579_ rbzero.wall_tracer.rayAddendY\[7\] _08447_ _01865_ _01714_ vssd1 vssd1 vccd1
+ vccd1 _01866_ sky130_fd_sc_hd__a22o_1
XFILLER_91_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19318_ rbzero.traced_texa\[-1\] rbzero.texV\[-1\] vssd1 vssd1 vccd1 vccd1 _02805_
+ sky130_fd_sc_hd__nor2_1
XFILLER_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09904_ rbzero.tex_r0\[46\] rbzero.tex_r0\[45\] _02995_ vssd1 vssd1 vccd1 vccd1 _03004_
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20024_ clknet_leaf_87_i_clk _00955_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09835_ _02966_ vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09766_ rbzero.tex_r1\[45\] rbzero.tex_r1\[46\] _02921_ vssd1 vssd1 vccd1 vccd1 _02930_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _03395_ _03343_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__or2_1
XFILLER_23_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11590_ rbzero.tex_b0\[13\] rbzero.tex_b0\[12\] _03732_ vssd1 vssd1 vccd1 vccd1 _04372_
+ sky130_fd_sc_hd__mux2_1
XFILLER_195_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10541_ _03337_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__buf_6
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13260_ _05469_ _06007_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__nor2_1
XFILLER_194_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10472_ _03143_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__clkbuf_4
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12211_ rbzero.wall_tracer.trackDistY\[-7\] vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__inv_2
XFILLER_170_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13191_ _05944_ _05947_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__xnor2_1
XFILLER_108_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12142_ _04855_ _04903_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__xor2_2
XFILLER_68_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16950_ _09553_ _09554_ vssd1 vssd1 vccd1 vccd1 _09556_ sky130_fd_sc_hd__nand2_1
X_12073_ _04837_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15901_ _03341_ vssd1 vssd1 vccd1 vccd1 _08524_ sky130_fd_sc_hd__clkbuf_4
X_11024_ rbzero.row_render.size\[0\] _03527_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__or2_1
X_16881_ _09486_ _09487_ vssd1 vssd1 vccd1 vccd1 _09488_ sky130_fd_sc_hd__nor2_1
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18620_ _02529_ vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__clkbuf_1
X_15832_ rbzero.wall_tracer.state\[14\] _03484_ _08450_ vssd1 vssd1 vccd1 vccd1 _08464_
+ sky130_fd_sc_hd__nand3_4
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18551_ rbzero.pov.spi_buffer\[44\] rbzero.pov.spi_buffer\[45\] _02488_ vssd1 vssd1
+ vccd1 vccd1 _02494_ sky130_fd_sc_hd__mux2_1
X_15763_ _08442_ vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__clkbuf_1
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ _05731_ _05528_ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__and2b_1
XFILLER_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17502_ _01790_ _01793_ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__xnor2_1
X_14714_ _07000_ _07401_ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__xnor2_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18482_ rbzero.pov.spi_buffer\[11\] rbzero.pov.spi_buffer\[12\] _02455_ vssd1 vssd1
+ vccd1 vccd1 _02458_ sky130_fd_sc_hd__mux2_1
X_11926_ _04672_ _04314_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__nand2_1
X_15694_ _08357_ _08376_ vssd1 vssd1 vccd1 vccd1 _08377_ sky130_fd_sc_hd__xnor2_2
XFILLER_33_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _01726_ _01727_ _01729_ vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__o21ai_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _07332_ vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__clkbuf_4
XFILLER_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _04532_ _04632_ net48 vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__a21o_1
XFILLER_60_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10808_ _03563_ _03567_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__nor2_1
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17364_ _01674_ vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14576_ _06857_ _06875_ _07007_ _07049_ vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__or4_1
XFILLER_60_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11788_ net18 _04564_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__nor2_1
X_16315_ _08807_ _08926_ vssd1 vssd1 vccd1 vccd1 _08927_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13527_ _06281_ _06283_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__nand2_1
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10739_ _03523_ _03524_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__or2_1
X_17295_ rbzero.wall_tracer.trackDistY\[5\] rbzero.wall_tracer.stepDistY\[5\] vssd1
+ vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__nor2_1
XFILLER_186_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16246_ _08856_ _08857_ vssd1 vssd1 vccd1 vccd1 _08858_ sky130_fd_sc_hd__nor2_1
XFILLER_158_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13458_ _06212_ _06214_ vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__nor2_1
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12409_ _05155_ _05156_ _05161_ _05163_ _05165_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__o2111a_1
X_16177_ _08245_ _08134_ _08260_ _08247_ vssd1 vssd1 vccd1 vccd1 _08790_ sky130_fd_sc_hd__o22a_1
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13389_ _06099_ _06143_ _06144_ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__a21oi_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15128_ rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerX\[-8\] _06850_
+ vssd1 vssd1 vccd1 vccd1 _07816_ sky130_fd_sc_hd__mux2_1
XFILLER_173_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19936_ net165 _00867_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[16\] sky130_fd_sc_hd__dfxtp_1
X_15059_ _07158_ _07167_ vssd1 vssd1 vccd1 vccd1 _07747_ sky130_fd_sc_hd__or2_1
XFILLER_123_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19867_ clknet_leaf_25_i_clk _00798_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_110_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18818_ rbzero.pov.ready_buffer\[13\] _02663_ _02670_ _02643_ vssd1 vssd1 vccd1 vccd1
+ _01050_ sky130_fd_sc_hd__o211a_1
XFILLER_95_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19798_ clknet_leaf_17_i_clk _00729_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_18405__47 clknet_1_0__leaf__02436_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__inv_2
XFILLER_83_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18749_ _02625_ _02627_ _02266_ vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__o21a_1
XFILLER_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_opt_1_0_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_1_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_192_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18914__100 clknet_1_1__leaf__02723_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__inv_2
XFILLER_132_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20007_ clknet_leaf_75_i_clk _00938_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_09818_ _02957_ vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__clkbuf_1
XFILLER_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09749_ _02909_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__clkbuf_4
XFILLER_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12760_ _05355_ _05469_ _05235_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__o21ai_4
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _04487_ net67 _04488_ net7 vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__a211o_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _05116_ _05447_ _05349_ _05310_ _05381_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__a32o_2
XFILLER_70_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _06893_ _07117_ vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__or2_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11642_ _03689_ _04418_ _04422_ _03679_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__a211o_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18960__142 clknet_1_1__leaf__02727_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__inv_2
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14361_ _07048_ vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__clkbuf_4
XFILLER_195_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11573_ rbzero.tex_b0\[21\] rbzero.tex_b0\[20\] _04189_ vssd1 vssd1 vccd1 vccd1 _04355_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16100_ _08294_ _08297_ vssd1 vssd1 vccd1 vccd1 _08714_ sky130_fd_sc_hd__nand2_1
Xinput18 i_gpout2_sel[3] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_6
XFILLER_11_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13312_ _05901_ _05904_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__and2_1
X_17080_ _09683_ _09684_ vssd1 vssd1 vccd1 vccd1 _09685_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10524_ _03329_ vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__clkbuf_1
Xinput29 i_gpout4_sel[2] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__buf_6
XFILLER_7_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14292_ rbzero.debug_overlay.playerY\[-3\] _06956_ vssd1 vssd1 vccd1 vccd1 _06980_
+ sky130_fd_sc_hd__or2_1
XFILLER_183_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16031_ _08642_ _08644_ vssd1 vssd1 vccd1 vccd1 _08645_ sky130_fd_sc_hd__and2_1
X_19056__228 clknet_1_1__leaf__02737_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__inv_2
X_13243_ _05997_ _05999_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__or2_1
X_10455_ _03293_ vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13174_ _05878_ _05880_ _05929_ _05930_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__o22ai_1
XFILLER_163_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10386_ _03257_ vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12125_ _04865_ _04869_ _04872_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__and3_1
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17982_ rbzero.pov.spi_buffer\[44\] rbzero.pov.ready_buffer\[44\] _02186_ vssd1 vssd1
+ vccd1 vccd1 _02192_ sky130_fd_sc_hd__mux2_1
X_19721_ clknet_leaf_87_i_clk _00652_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16933_ _09468_ _09538_ vssd1 vssd1 vccd1 vccd1 _09539_ sky130_fd_sc_hd__nand2_1
XFILLER_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12056_ _02907_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__buf_4
XFILLER_46_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11007_ rbzero.row_render.size\[9\] _03778_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__nor2_1
XFILLER_77_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19652_ clknet_leaf_18_i_clk _00583_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16864_ _09465_ _09470_ vssd1 vssd1 vccd1 vccd1 _09471_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18603_ rbzero.pov.spi_buffer\[69\] rbzero.pov.spi_buffer\[70\] _02443_ vssd1 vssd1
+ vccd1 vccd1 _02521_ sky130_fd_sc_hd__mux2_1
X_15815_ rbzero.traced_texa\[-4\] _08461_ _08459_ rbzero.wall_tracer.visualWallDist\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__a22o_1
X_16795_ _09208_ _09402_ vssd1 vssd1 vccd1 vccd1 _09403_ sky130_fd_sc_hd__nand2_1
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19583_ clknet_leaf_61_i_clk _00514_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15746_ _08427_ _08428_ vssd1 vssd1 vccd1 vccd1 _08429_ sky130_fd_sc_hd__nor2_2
X_18534_ rbzero.pov.spi_buffer\[36\] rbzero.pov.spi_buffer\[37\] _02477_ vssd1 vssd1
+ vccd1 vccd1 _02485_ sky130_fd_sc_hd__mux2_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ _05701_ _05712_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__and2b_1
XFILLER_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11909_ _04532_ _04666_ _04668_ net53 _04683_ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__a221o_1
X_15677_ _07281_ _08000_ _07123_ _06858_ vssd1 vssd1 vccd1 vccd1 _08360_ sky130_fd_sc_hd__o22a_1
X_18465_ rbzero.pov.spi_buffer\[3\] rbzero.pov.spi_buffer\[4\] _02444_ vssd1 vssd1
+ vccd1 vccd1 _02449_ sky130_fd_sc_hd__mux2_1
X_12889_ _05533_ _05645_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17416_ rbzero.debug_overlay.vplaneY\[-9\] _01714_ _08448_ rbzero.wall_tracer.rayAddendY\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__a22o_1
X_14628_ _07293_ _07307_ vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__and2b_1
XFILLER_178_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17347_ rbzero.spi_registers.new_mapd\[2\] rbzero.spi_registers.spi_buffer\[2\] _01663_
+ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__mux2_1
XFILLER_187_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14559_ _06969_ _07024_ vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__or2_1
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17278_ _01534_ _01605_ _01607_ _01526_ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__a31o_1
XFILLER_146_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16229_ rbzero.wall_tracer.trackDistX\[1\] _08553_ _08835_ _08841_ vssd1 vssd1 vccd1
+ vccd1 _00550_ sky130_fd_sc_hd__o22a_1
XFILLER_127_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19919_ clknet_leaf_96_i_clk _00850_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19161__323 clknet_1_0__leaf__02747_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__inv_2
XFILLER_58_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20487_ clknet_leaf_40_i_clk _01418_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10240_ rbzero.tex_g0\[15\] rbzero.tex_g0\[14\] _03177_ vssd1 vssd1 vccd1 vccd1 _03181_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10171_ rbzero.tex_g0\[48\] rbzero.tex_g0\[47\] _03144_ vssd1 vssd1 vccd1 vccd1 _03145_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13930_ _05271_ _06636_ _06681_ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__o21a_1
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13861_ _06601_ _06617_ vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__nor2_1
X_15600_ _08243_ _08283_ vssd1 vssd1 vccd1 vccd1 _08284_ sky130_fd_sc_hd__nand2_1
XFILLER_41_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12812_ _05556_ _05566_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__or2_1
XFILLER_74_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16580_ _08970_ _09188_ vssd1 vssd1 vccd1 vccd1 _09190_ sky130_fd_sc_hd__or2_1
X_13792_ _06539_ _06548_ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__nand2_1
XFILLER_76_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15531_ _08075_ _08086_ _08084_ vssd1 vssd1 vccd1 vccd1 _08215_ sky130_fd_sc_hd__a21oi_1
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12743_ _05492_ _05497_ _05498_ _05499_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__a22o_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18250_ rbzero.spi_registers.vshift\[4\] _02349_ vssd1 vssd1 vccd1 vccd1 _02354_
+ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_91_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15462_ _08138_ _08143_ _08146_ vssd1 vssd1 vccd1 vccd1 _08147_ sky130_fd_sc_hd__and3_1
XFILLER_176_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12674_ _05414_ _05346_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__or2_1
XFILLER_30_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ rbzero.wall_tracer.trackDistY\[-8\] rbzero.wall_tracer.stepDistY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__or2_1
X_14413_ _06917_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__buf_2
XFILLER_179_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11625_ _04192_ _04403_ _04405_ _04179_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__o211a_1
X_18181_ rbzero.spi_registers.new_mapd\[0\] _02289_ _02308_ _02301_ vssd1 vssd1 vccd1
+ vccd1 _00775_ sky130_fd_sc_hd__o211a_1
X_15393_ _06979_ _07332_ vssd1 vssd1 vccd1 vccd1 _08078_ sky130_fd_sc_hd__nor2_1
XFILLER_168_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17132_ _09632_ _09656_ _01475_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__a21oi_1
XFILLER_184_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14344_ rbzero.debug_overlay.playerX\[-1\] rbzero.debug_overlay.playerX\[-2\] _06987_
+ vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__or3_4
X_11556_ rbzero.tex_b0\[37\] rbzero.tex_b0\[36\] _04189_ vssd1 vssd1 vccd1 vccd1 _04338_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17063_ _09666_ _09667_ vssd1 vssd1 vccd1 vccd1 _09668_ sky130_fd_sc_hd__nor2_1
X_10507_ _03320_ vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14275_ _06961_ _06962_ vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__nand2_1
X_11487_ rbzero.tex_g1\[1\] rbzero.tex_g1\[0\] _03727_ vssd1 vssd1 vccd1 vccd1 _04270_
+ sky130_fd_sc_hd__mux2_1
XFILLER_144_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16014_ _08336_ _08345_ _08343_ vssd1 vssd1 vccd1 vccd1 _08628_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_0__02752_ _02752_ vssd1 vssd1 vccd1 vccd1 clknet_0__02752_ sky130_fd_sc_hd__clkbuf_16
X_13226_ _05945_ _05944_ _05981_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__a21oi_1
X_10438_ _03284_ vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13157_ _05355_ _05503_ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__nor2_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _03248_ vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__clkbuf_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12108_ rbzero.debug_overlay.facingY\[-1\] rbzero.wall_tracer.rayAddendY\[7\] vssd1
+ vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__and2_1
XFILLER_112_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _05831_ _05825_ _05829_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__or3_1
X_17965_ rbzero.pov.spi_buffer\[36\] rbzero.pov.ready_buffer\[36\] _02175_ vssd1 vssd1
+ vccd1 vccd1 _02183_ sky130_fd_sc_hd__mux2_1
XFILLER_2_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19704_ clknet_leaf_71_i_clk _00635_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12039_ _03838_ _02901_ _04779_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__mux2_1
X_16916_ _09521_ _09522_ vssd1 vssd1 vccd1 vccd1 _09523_ sky130_fd_sc_hd__and2b_1
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17896_ rbzero.pov.spi_buffer\[3\] rbzero.pov.ready_buffer\[3\] _02143_ vssd1 vssd1
+ vccd1 vccd1 _02147_ sky130_fd_sc_hd__mux2_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19110__277 clknet_1_0__leaf__02742_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_44_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19635_ clknet_leaf_59_i_clk _00566_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16847_ _09452_ _09453_ vssd1 vssd1 vccd1 vccd1 _09454_ sky130_fd_sc_hd__or2_1
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18967__148 clknet_1_1__leaf__02728_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__inv_2
XFILLER_19_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19566_ clknet_leaf_35_i_clk _00497_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16778_ _09283_ _09385_ vssd1 vssd1 vccd1 vccd1 _09386_ sky130_fd_sc_hd__xnor2_1
XFILLER_168_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18517_ rbzero.pov.spi_buffer\[28\] rbzero.pov.spi_buffer\[29\] _02466_ vssd1 vssd1
+ vccd1 vccd1 _02476_ sky130_fd_sc_hd__mux2_1
X_15729_ _08258_ _08280_ _08278_ vssd1 vssd1 vccd1 vccd1 _08412_ sky130_fd_sc_hd__a21oi_1
XFILLER_178_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19497_ clknet_leaf_47_i_clk _00443_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_179_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_59_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18448_ clknet_1_0__leaf__04486_ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__buf_1
XFILLER_61_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18379_ _02421_ _02430_ _02431_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__and3_1
XFILLER_30_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20410_ net470 _01341_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19004__182 clknet_1_0__leaf__02731_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__inv_2
XFILLER_175_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20341_ net401 _01272_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20272_ net332 _01203_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__02741_ clknet_0__02741_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02741_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_99_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11410_ rbzero.tex_g0\[51\] _03729_ _03730_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__and3_1
XFILLER_165_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12390_ _05138_ _05140_ _05146_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__a21o_1
XFILLER_193_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_74 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_74/HI o_rgb[1] sky130_fd_sc_hd__conb_1
XFILLER_193_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_85 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_85/HI o_rgb[16] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_96 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_96/HI zeros[5] sky130_fd_sc_hd__conb_1
XFILLER_181_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11341_ rbzero.debug_overlay.playerX\[5\] _04125_ _03519_ gpout0.vpos\[3\] vssd1
+ vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__a211o_1
XFILLER_180_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14060_ rbzero.wall_tracer.trackDistY\[-9\] _06786_ _06792_ vssd1 vssd1 vccd1 vccd1
+ _00430_ sky130_fd_sc_hd__o21a_1
X_11272_ gpout0.hpos\[4\] _04040_ _04052_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__or3_1
XFILLER_152_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13011_ _05467_ _05483_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__nand2_2
X_10223_ rbzero.tex_g0\[23\] rbzero.tex_g0\[22\] _03166_ vssd1 vssd1 vccd1 vccd1 _03172_
+ sky130_fd_sc_hd__mux2_1
X_19248__22 clknet_1_0__leaf__02755_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__inv_2
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10154_ _03135_ vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19168__329 clknet_1_1__leaf__02748_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__inv_2
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14962_ _07621_ _07649_ vssd1 vssd1 vccd1 vccd1 _07650_ sky130_fd_sc_hd__xnor2_1
X_17750_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.debug_overlay.vplaneX\[-6\] _02016_
+ _02017_ vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10085_ _03099_ vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16701_ rbzero.wall_tracer.trackDistX\[5\] rbzero.wall_tracer.stepDistX\[5\] vssd1
+ vssd1 vccd1 vccd1 _09310_ sky130_fd_sc_hd__and2_1
XFILLER_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13913_ _05376_ _06666_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__nor2_1
X_14893_ _06968_ vssd1 vssd1 vccd1 vccd1 _07581_ sky130_fd_sc_hd__buf_2
X_17681_ _01951_ _01952_ _01954_ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__or3_1
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19420_ _01703_ _01711_ _01710_ _08464_ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__a31o_1
X_16632_ _09111_ _09120_ _09118_ vssd1 vssd1 vccd1 vccd1 _09241_ sky130_fd_sc_hd__a21oi_1
X_13844_ _05349_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__buf_2
XFILLER_62_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19351_ _02759_ _02832_ _02833_ _02319_ rbzero.texV\[3\] vssd1 vssd1 vccd1 vccd1
+ _01420_ sky130_fd_sc_hd__a32o_1
X_16563_ _09045_ _09057_ _09055_ vssd1 vssd1 vccd1 vccd1 _09173_ sky130_fd_sc_hd__a21oi_2
X_13775_ _06122_ _06230_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__or2_1
X_10987_ rbzero.row_render.size\[3\] _03772_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__or2_1
XFILLER_31_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18302_ _02384_ vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__clkbuf_1
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15514_ _08192_ _08197_ vssd1 vssd1 vccd1 vccd1 _08198_ sky130_fd_sc_hd__xnor2_1
X_12726_ _05482_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__clkbuf_2
X_16494_ _09102_ _09103_ vssd1 vssd1 vccd1 vccd1 _09104_ sky130_fd_sc_hd__nor2_1
XFILLER_31_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19282_ _02774_ _02775_ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__xnor2_1
XFILLER_71_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15445_ _07748_ vssd1 vssd1 vccd1 vccd1 _08130_ sky130_fd_sc_hd__buf_2
X_18233_ _02343_ vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__clkbuf_1
X_12657_ _05269_ _05320_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__nand2_2
XFILLER_129_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11608_ _04018_ _04028_ _04311_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__o21a_1
XFILLER_157_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15376_ _07940_ _08047_ vssd1 vssd1 vccd1 vccd1 _08061_ sky130_fd_sc_hd__nor2_1
X_18164_ rbzero.spi_registers.new_mapd\[4\] _02290_ _02299_ _02275_ vssd1 vssd1 vccd1
+ vccd1 _00767_ sky130_fd_sc_hd__o211a_1
XFILLER_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12588_ _05197_ _05257_ _05313_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__mux2_1
XFILLER_11_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17115_ _09693_ _09698_ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__or2b_1
X_14327_ _06876_ _07014_ vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__nand2_1
XFILLER_156_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11539_ rbzero.tex_b0\[61\] rbzero.tex_b0\[60\] _04189_ vssd1 vssd1 vccd1 vccd1 _04321_
+ sky130_fd_sc_hd__mux2_1
X_18095_ _02252_ vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17046_ _09635_ _09650_ vssd1 vssd1 vccd1 vccd1 _09651_ sky130_fd_sc_hd__and2_1
X_14258_ rbzero.debug_overlay.playerX\[-5\] _06927_ vssd1 vssd1 vccd1 vccd1 _06946_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_172_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__02735_ _02735_ vssd1 vssd1 vccd1 vccd1 clknet_0__02735_ sky130_fd_sc_hd__clkbuf_16
X_13209_ _05928_ _05963_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__and2_1
XFILLER_171_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ rbzero.debug_overlay.playerY\[-7\] rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerY\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__or3_1
XFILLER_97_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18447__86 clknet_1_0__leaf__02439_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__inv_2
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ rbzero.pov.spi_buffer\[28\] rbzero.pov.ready_buffer\[28\] _02164_ vssd1 vssd1
+ vccd1 vccd1 _02174_ sky130_fd_sc_hd__mux2_1
XFILLER_100_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17879_ rbzero.spi_registers.spi_counter\[4\] _02102_ _02103_ _02135_ vssd1 vssd1
+ vccd1 vccd1 _00646_ sky130_fd_sc_hd__o211a_1
XFILLER_94_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19618_ clknet_leaf_47_i_clk _00549_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_199_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19549_ clknet_leaf_33_i_clk _00480_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20324_ net384 _01255_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20255_ net315 _01186_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20186_ net246 _01117_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09997_ rbzero.tex_r0\[2\] rbzero.tex_r0\[1\] _03050_ vssd1 vssd1 vccd1 vccd1 _03053_
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10910_ _03556_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__buf_4
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11890_ net22 net21 vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__and2b_1
Xclkbuf_1_0__f__02724_ clknet_0__02724_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02724_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10841_ _03595_ _03603_ _03622_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__nor3_4
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13560_ _06173_ _06315_ _06316_ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__a21bo_1
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10772_ _03556_ _03557_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__nor2_2
XFILLER_71_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12511_ _05235_ _05244_ _05267_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__and3_1
XFILLER_73_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13491_ _06148_ _06247_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15230_ _07914_ _07915_ vssd1 vssd1 vccd1 vccd1 _07917_ sky130_fd_sc_hd__nand2_1
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12442_ _05187_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__buf_2
XFILLER_60_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15161_ _07724_ _07833_ _07846_ vssd1 vssd1 vccd1 vccd1 _07848_ sky130_fd_sc_hd__and3_1
XFILLER_126_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12373_ rbzero.wall_tracer.rcp_sel\[2\] _04899_ _04900_ vssd1 vssd1 vccd1 vccd1 _05130_
+ sky130_fd_sc_hd__and3_1
XFILLER_197_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14112_ _06820_ vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__clkbuf_1
X_11324_ rbzero.debug_overlay.vplaneY\[-2\] vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__clkbuf_4
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15092_ _07778_ _07779_ vssd1 vssd1 vccd1 vccd1 _07780_ sky130_fd_sc_hd__nor2_2
XFILLER_107_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14043_ rbzero.wall_tracer.stepDistY\[9\] _06779_ _04836_ vssd1 vssd1 vccd1 vccd1
+ _06780_ sky130_fd_sc_hd__mux2_1
XFILLER_10_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11255_ _04039_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__buf_2
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10206_ rbzero.tex_g0\[31\] rbzero.tex_g0\[30\] _03155_ vssd1 vssd1 vccd1 vccd1 _03163_
+ sky130_fd_sc_hd__mux2_1
XFILLER_140_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18851_ _04109_ _02634_ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__and2_1
XFILLER_80_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11186_ rbzero.tex_r1\[12\] _03920_ _03925_ _03969_ _03970_ vssd1 vssd1 vccd1 vccd1
+ _03971_ sky130_fd_sc_hd__a311o_1
XFILLER_192_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17802_ _02064_ _02065_ _02062_ _02063_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__o211ai_2
XFILLER_67_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10137_ _03126_ vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__clkbuf_1
X_18782_ _03338_ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__clkbuf_4
X_15994_ _07856_ _08070_ vssd1 vssd1 vccd1 vccd1 _08608_ sky130_fd_sc_hd__nor2_1
XFILLER_0_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17733_ _01986_ _01990_ _02002_ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__a21oi_1
X_14945_ _07541_ _07632_ vssd1 vssd1 vccd1 vccd1 _07633_ sky130_fd_sc_hd__xor2_1
X_10068_ _03090_ vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17664_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.debug_overlay.vplaneX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__nand2_1
XFILLER_36_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14876_ _07548_ _07563_ vssd1 vssd1 vccd1 vccd1 _07564_ sky130_fd_sc_hd__nor2_1
X_19403_ rbzero.traced_texVinit\[9\] _02868_ _08454_ _08834_ vssd1 vssd1 vccd1 vccd1
+ _01437_ sky130_fd_sc_hd__a22o_1
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16615_ _09222_ _09223_ vssd1 vssd1 vccd1 vccd1 _09224_ sky130_fd_sc_hd__nor2_1
XFILLER_78_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13827_ _06224_ _06583_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__and2_1
X_17595_ _01786_ rbzero.wall_tracer.rayAddendY\[9\] vssd1 vssd1 vccd1 vccd1 _01880_
+ sky130_fd_sc_hd__or2_1
XFILLER_189_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19334_ _02816_ _02817_ _02818_ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__and3_1
X_16546_ _08247_ _08245_ _09036_ _08678_ vssd1 vssd1 vccd1 vccd1 _09156_ sky130_fd_sc_hd__nor4_1
X_13758_ _06337_ _06513_ vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__nand2_1
XFILLER_43_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19222__378 clknet_1_0__leaf__02753_ vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__inv_2
XFILLER_189_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12709_ _05450_ _05458_ _05465_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__a21bo_1
X_19265_ _03338_ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__buf_4
X_13689_ _06440_ _06443_ _06445_ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__a21oi_1
X_16477_ _08562_ _09086_ _09087_ _08487_ vssd1 vssd1 vccd1 vccd1 _09088_ sky130_fd_sc_hd__a31o_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18216_ _02331_ vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__clkbuf_1
X_15428_ _08101_ _08112_ vssd1 vssd1 vccd1 vccd1 _08113_ sky130_fd_sc_hd__xor2_1
XFILLER_15_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15359_ _07941_ _08044_ vssd1 vssd1 vccd1 vccd1 _08045_ sky130_fd_sc_hd__xnor2_4
X_18147_ rbzero.spi_registers.got_new_mapd _02288_ vssd1 vssd1 vccd1 vccd1 _02289_
+ sky130_fd_sc_hd__nand2_2
XFILLER_156_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18078_ rbzero.spi_registers.spi_buffer\[15\] rbzero.spi_registers.spi_buffer\[14\]
+ _02226_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__mux2_1
XFILLER_172_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09920_ _03012_ vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17029_ _09534_ vssd1 vssd1 vccd1 vccd1 _09634_ sky130_fd_sc_hd__inv_2
XFILLER_172_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20040_ clknet_leaf_5_i_clk _00971_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_19116__283 clknet_1_1__leaf__02742_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__inv_2
X_09851_ _02974_ vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__clkbuf_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09782_ _02938_ vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__clkbuf_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__02440_ clknet_0__02440_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02440_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_139_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20307_ net367 _01238_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11040_ rbzero.floor_leak\[3\] _03624_ _03673_ rbzero.floor_leak\[2\] _03825_ vssd1
+ vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__o221a_1
XFILLER_89_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20238_ net298 _01169_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20169_ net229 _01100_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _05729_ _05747_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__xnor2_1
XFILLER_58_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14730_ _07072_ _07417_ vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__nand2_1
X_11942_ net44 _04665_ _04685_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__and3_1
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _07296_ _07344_ _07345_ _07348_ vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__o2bb2a_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _03459_ _03469_ _04612_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__mux2_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16400_ _08885_ _09008_ _09010_ vssd1 vssd1 vccd1 vccd1 _09011_ sky130_fd_sc_hd__a21bo_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ _06122_ _05987_ _06368_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__o21ba_1
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10824_ _03609_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__buf_4
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14592_ _07278_ _07279_ vssd1 vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__or2_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17380_ _08509_ _08473_ _01682_ _01683_ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__a31o_1
XFILLER_60_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16331_ _08882_ _08942_ vssd1 vssd1 vccd1 vccd1 _08943_ sky130_fd_sc_hd__xnor2_1
X_13543_ _06247_ _06296_ _06299_ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__a21o_1
X_10755_ _03538_ _03540_ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__nand2_1
XFILLER_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16262_ _08861_ _08873_ vssd1 vssd1 vccd1 vccd1 _08874_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13474_ _05472_ _06230_ vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__or2_1
XFILLER_186_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10686_ _03478_ _03340_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__nor2_1
XFILLER_199_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15213_ _07185_ _07897_ vssd1 vssd1 vccd1 vccd1 _07900_ sky130_fd_sc_hd__nor2_1
X_18001_ rbzero.pov.spi_buffer\[53\] rbzero.pov.ready_buffer\[53\] _02197_ vssd1 vssd1
+ vccd1 vccd1 _02202_ sky130_fd_sc_hd__mux2_1
X_12425_ _05178_ _05180_ _05181_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__and3b_1
XFILLER_200_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16193_ _08804_ _08805_ vssd1 vssd1 vccd1 vccd1 _08806_ sky130_fd_sc_hd__and2b_1
XFILLER_138_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15144_ _07805_ _07806_ vssd1 vssd1 vccd1 vccd1 _07831_ sky130_fd_sc_hd__and2b_1
XFILLER_127_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12356_ _05040_ _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__and2_1
XFILLER_181_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ _04051_ _04091_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__nor2_4
X_19952_ net181 _00883_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[32\] sky130_fd_sc_hd__dfxtp_1
X_15075_ _07760_ _07762_ vssd1 vssd1 vccd1 vccd1 _07763_ sky130_fd_sc_hd__xor2_2
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12287_ _05040_ _05041_ _05042_ _05043_ vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__o211a_1
X_18903_ rbzero.spi_registers.got_new_mapd _02323_ _02283_ _01663_ vssd1 vssd1 vccd1
+ vccd1 _01083_ sky130_fd_sc_hd__a31o_1
X_14026_ _06766_ vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11238_ gpout0.vpos\[6\] _03460_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__xnor2_1
X_19883_ clknet_leaf_22_i_clk _00814_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18834_ rbzero.pov.ready_buffer\[20\] _02663_ _02679_ _02672_ vssd1 vssd1 vccd1 vccd1
+ _01057_ sky130_fd_sc_hd__o211a_1
XFILLER_171_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11169_ rbzero.tex_r1\[33\] _03659_ _03767_ _03634_ vssd1 vssd1 vccd1 vccd1 _03954_
+ sky130_fd_sc_hd__a31o_1
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__02434_ _02434_ vssd1 vssd1 vccd1 vccd1 clknet_0__02434_ sky130_fd_sc_hd__clkbuf_16
XFILLER_83_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18765_ rbzero.pov.ready_buffer\[34\] _02636_ _02640_ _02586_ vssd1 vssd1 vccd1 vccd1
+ _01027_ sky130_fd_sc_hd__o211a_1
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15977_ rbzero.wall_tracer.trackDistX\[-1\] _08553_ _08585_ _08591_ vssd1 vssd1 vccd1
+ vccd1 _00548_ sky130_fd_sc_hd__o22a_1
XFILLER_49_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17716_ rbzero.debug_overlay.vplaneX\[10\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__or2_1
X_14928_ _06866_ _07100_ vssd1 vssd1 vccd1 vccd1 _07616_ sky130_fd_sc_hd__or2_1
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18696_ net40 _02532_ _02262_ vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__o21a_2
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17647_ _01922_ _01923_ vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__nand2_1
X_14859_ _07544_ _07546_ vssd1 vssd1 vccd1 vccd1 _07547_ sky130_fd_sc_hd__nor2_1
XFILLER_63_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17578_ _01863_ _01864_ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__xor2_1
X_19317_ _02759_ _02803_ _02804_ _02319_ rbzero.texV\[-2\] vssd1 vssd1 vccd1 vccd1
+ _01415_ sky130_fd_sc_hd__a32o_1
XFILLER_91_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16529_ _09014_ _09016_ _08134_ _08260_ vssd1 vssd1 vccd1 vccd1 _09139_ sky130_fd_sc_hd__or4_1
XFILLER_149_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09903_ _03003_ vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09834_ rbzero.tex_r1\[13\] rbzero.tex_r1\[14\] _02965_ vssd1 vssd1 vccd1 vccd1 _02966_
+ sky130_fd_sc_hd__mux2_1
X_20023_ clknet_leaf_88_i_clk _00954_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09765_ _02929_ vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10540_ _02981_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__buf_4
XFILLER_168_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10471_ _03301_ vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__clkbuf_1
XFILLER_157_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12210_ rbzero.wall_tracer.trackDistY\[-6\] vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__inv_2
XFILLER_182_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13190_ _05945_ _05946_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__nor2_1
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12141_ _04857_ _04864_ _04852_ _04850_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__a31o_1
XFILLER_2_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12072_ net72 rbzero.wall_tracer.state\[12\] _04834_ vssd1 vssd1 vccd1 vccd1 _04837_
+ sky130_fd_sc_hd__and3_1
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11023_ gpout0.hpos\[1\] gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__or2_1
X_15900_ rbzero.wall_tracer.trackDistX\[-10\] _08508_ _08517_ _08523_ vssd1 vssd1
+ vccd1 vccd1 _00539_ sky130_fd_sc_hd__o22a_1
X_16880_ _09016_ _09036_ _09046_ _09014_ vssd1 vssd1 vccd1 vccd1 _09487_ sky130_fd_sc_hd__o22a_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15831_ rbzero.traced_texa\[10\] _08463_ _08462_ rbzero.wall_tracer.visualWallDist\[10\]
+ vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__a22o_1
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18550_ _02493_ vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ _05495_ _05727_ _05730_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__o21a_1
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15762_ _03502_ _08441_ _08439_ vssd1 vssd1 vccd1 vccd1 _08442_ sky130_fd_sc_hd__and3_1
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ _01791_ _01779_ _01792_ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__a21o_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14713_ _06993_ _07005_ vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__nor2_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18481_ _02457_ vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11925_ _04677_ _04681_ _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__o21ai_2
X_15693_ _08358_ _08375_ vssd1 vssd1 vccd1 vccd1 _08376_ sky130_fd_sc_hd__xor2_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _01728_ _01718_ _01717_ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__a21oi_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14644_ rbzero.wall_tracer.visualWallDist\[4\] _06855_ vssd1 vssd1 vccd1 vccd1 _07332_
+ sky130_fd_sc_hd__nand2_2
X_11856_ net14 net13 vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__nor2_1
XFILLER_127_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10807_ _03591_ _03592_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__xnor2_1
X_14575_ _07237_ _07241_ vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__or2b_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17363_ rbzero.spi_registers.new_mapd\[10\] rbzero.spi_registers.spi_buffer\[10\]
+ _01662_ vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__mux2_1
X_11787_ net17 vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__inv_2
XFILLER_41_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16314_ _08923_ _08925_ vssd1 vssd1 vccd1 vccd1 _08926_ sky130_fd_sc_hd__xor2_1
XFILLER_174_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10738_ gpout0.hpos\[4\] vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__clkbuf_4
X_13526_ _06211_ _06282_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__or2_1
X_17294_ rbzero.wall_tracer.trackDistY\[4\] _01558_ _01621_ _09197_ vssd1 vssd1 vccd1
+ vccd1 _00575_ sky130_fd_sc_hd__o22a_1
X_16245_ _08854_ _08855_ vssd1 vssd1 vccd1 vccd1 _08857_ sky130_fd_sc_hd__and2_1
XFILLER_146_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13457_ _06196_ _06213_ vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__nor2_1
X_10669_ _03463_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__buf_4
XFILLER_127_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12408_ _05164_ _05067_ _03489_ _05078_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__a211o_1
XFILLER_126_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16176_ _08245_ _08260_ _08380_ vssd1 vssd1 vccd1 vccd1 _08789_ sky130_fd_sc_hd__nor3_1
XFILLER_154_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13388_ _06099_ _06143_ _06144_ vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__and3_1
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12339_ _05034_ _05095_ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__xnor2_2
X_15127_ _07699_ _07528_ vssd1 vssd1 vccd1 vccd1 _07815_ sky130_fd_sc_hd__xor2_4
XFILLER_126_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19033__207 clknet_1_1__leaf__02735_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__inv_2
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19935_ net164 _00866_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[15\] sky130_fd_sc_hd__dfxtp_1
X_15058_ _07744_ _07745_ vssd1 vssd1 vccd1 vccd1 _07746_ sky130_fd_sc_hd__xnor2_2
XFILLER_130_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14009_ _05476_ _06749_ _06751_ _05373_ _06693_ vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__a32o_1
X_19866_ clknet_leaf_24_i_clk _00797_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18817_ rbzero.debug_overlay.vplaneX\[-7\] _02660_ vssd1 vssd1 vccd1 vccd1 _02670_
+ sky130_fd_sc_hd__or2_1
XFILLER_23_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19797_ clknet_leaf_17_i_clk _00728_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_23_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18748_ rbzero.pov.ready_buffer\[57\] _02540_ _02588_ _02626_ vssd1 vssd1 vccd1 vccd1
+ _02627_ sky130_fd_sc_hd__o211a_1
XFILLER_23_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19228__384 clknet_1_0__leaf__02753_ vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__inv_2
XFILLER_37_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18679_ rbzero.debug_overlay.playerX\[3\] _02533_ _02573_ _02559_ vssd1 vssd1 vccd1
+ vccd1 _01008_ sky130_fd_sc_hd__a211o_1
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20006_ clknet_leaf_75_i_clk _00937_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09817_ rbzero.tex_r1\[21\] rbzero.tex_r1\[22\] _02954_ vssd1 vssd1 vccd1 vccd1 _02957_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09748_ _02920_ vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _04487_ _03913_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__nor2_1
XFILLER_15_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12690_ _05270_ _05367_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__nor2_2
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _03693_ _04419_ _04420_ _04421_ _03673_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__o221a_1
XFILLER_39_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14360_ _07047_ vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__buf_2
X_11572_ rbzero.tex_b0\[23\] _04155_ _04156_ _03611_ vssd1 vssd1 vccd1 vccd1 _04354_
+ sky130_fd_sc_hd__a31o_1
XFILLER_161_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13311_ _05990_ _05995_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__nor2_1
XFILLER_168_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10523_ rbzero.tex_b0\[8\] rbzero.tex_b0\[7\] _03324_ vssd1 vssd1 vccd1 vccd1 _03329_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput19 i_gpout2_sel[4] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_8
XFILLER_196_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14291_ _06978_ vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__clkbuf_4
X_16030_ _08643_ _07857_ _08641_ vssd1 vssd1 vccd1 vccd1 _08644_ sky130_fd_sc_hd__o21ai_1
XFILLER_6_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13242_ _05993_ _05996_ _05998_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__a21oi_1
XFILLER_196_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10454_ rbzero.tex_b0\[41\] rbzero.tex_b0\[40\] _03291_ vssd1 vssd1 vccd1 vccd1 _03293_
+ sky130_fd_sc_hd__mux2_1
XFILLER_170_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13173_ _05493_ _05471_ _05926_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__o21a_1
X_10385_ rbzero.tex_b1\[9\] rbzero.tex_b1\[10\] _03254_ vssd1 vssd1 vccd1 vccd1 _03257_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12124_ _04884_ _04885_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__and2_1
XFILLER_2_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17981_ _02191_ vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19720_ clknet_leaf_95_i_clk _00651_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12055_ rbzero.hsync vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__inv_2
X_16932_ _09470_ _09465_ vssd1 vssd1 vccd1 vccd1 _09538_ sky130_fd_sc_hd__or2b_1
XFILLER_81_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11006_ _02900_ _03777_ _03780_ _02902_ _03791_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__a221o_1
X_19651_ clknet_leaf_16_i_clk _00582_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_mapd\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16863_ _09468_ _09469_ vssd1 vssd1 vccd1 vccd1 _09470_ sky130_fd_sc_hd__nand2_2
XFILLER_38_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18602_ _02520_ vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15814_ _08460_ vssd1 vssd1 vccd1 vccd1 _08461_ sky130_fd_sc_hd__clkbuf_4
XFILLER_65_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19582_ clknet_leaf_62_i_clk _00513_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16794_ _09400_ _09401_ vssd1 vssd1 vccd1 vccd1 _09402_ sky130_fd_sc_hd__xnor2_1
X_18533_ _02484_ vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15745_ _08424_ _08426_ vssd1 vssd1 vccd1 vccd1 _08428_ sky130_fd_sc_hd__and2_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _05693_ _05694_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__xnor2_1
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18464_ _02448_ vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11908_ net51 _04665_ _04669_ net50 vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__a22o_1
X_15676_ _06857_ _08000_ vssd1 vssd1 vccd1 vccd1 _08359_ sky130_fd_sc_hd__or2_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _05603_ _05644_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _03340_ vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__clkbuf_4
XFILLER_33_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14627_ _07309_ _07314_ vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11839_ _04612_ _04393_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__nor2_1
XFILLER_53_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17346_ _01665_ vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14558_ _07244_ _07245_ vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__nor2_1
XFILLER_53_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13509_ _06259_ _06264_ _06265_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__a21oi_1
XFILLER_174_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17277_ _01606_ vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__inv_2
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14489_ rbzero.wall_tracer.visualWallDist\[-10\] _06854_ vssd1 vssd1 vccd1 vccd1
+ _07177_ sky130_fd_sc_hd__nand2_2
XFILLER_174_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16228_ _08562_ _08839_ _08840_ _08522_ vssd1 vssd1 vccd1 vccd1 _08841_ sky130_fd_sc_hd__a31o_1
XFILLER_173_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16159_ _08770_ _08771_ vssd1 vssd1 vccd1 vccd1 _08772_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19918_ clknet_leaf_96_i_clk _00849_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19849_ clknet_leaf_24_i_clk _00780_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18944__127 clknet_1_0__leaf__02726_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__inv_2
XFILLER_145_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20486_ clknet_leaf_40_i_clk _01417_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10170_ _03143_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__clkbuf_4
XFILLER_117_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18990__169 clknet_1_1__leaf__02730_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__inv_2
XFILLER_78_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13860_ _06561_ _06616_ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12811_ _05499_ _05498_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__xnor2_1
X_13791_ _06531_ _06538_ vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__nand2_1
XFILLER_62_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18396__39 clknet_1_0__leaf__02435_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__inv_2
X_15530_ _08202_ _08213_ vssd1 vssd1 vccd1 vccd1 _08214_ sky130_fd_sc_hd__xnor2_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _05495_ _05433_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__nor2_2
XFILLER_16_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15461_ _07174_ _08144_ _08145_ vssd1 vssd1 vccd1 vccd1 _08146_ sky130_fd_sc_hd__a21o_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12673_ _05426_ _05429_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__nand2_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17200_ rbzero.wall_tracer.trackDistY\[-9\] _01523_ _01540_ _08525_ vssd1 vssd1 vccd1
+ vccd1 _00562_ sky130_fd_sc_hd__o22a_1
X_11624_ _03652_ _04404_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__or2_1
X_14412_ _06933_ vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__clkbuf_4
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18180_ rbzero.mapdyw\[0\] _02291_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__or2_1
X_15392_ _07856_ _07787_ vssd1 vssd1 vccd1 vccd1 _08077_ sky130_fd_sc_hd__nor2_1
XFILLER_156_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17131_ _09657_ _09690_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__and2b_1
XFILLER_168_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11555_ rbzero.tex_b0\[39\] _04155_ _04156_ _03611_ vssd1 vssd1 vccd1 vccd1 _04337_
+ sky130_fd_sc_hd__a31o_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14343_ rbzero.wall_tracer.visualWallDist\[-1\] _07030_ _03490_ vssd1 vssd1 vccd1
+ vccd1 _07031_ sky130_fd_sc_hd__mux2_1
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10506_ rbzero.tex_b0\[16\] rbzero.tex_b0\[15\] _03313_ vssd1 vssd1 vccd1 vccd1 _03320_
+ sky130_fd_sc_hd__mux2_1
X_17062_ _08888_ _08333_ _09568_ _09567_ vssd1 vssd1 vccd1 vccd1 _09667_ sky130_fd_sc_hd__o31a_1
X_14274_ rbzero.debug_overlay.playerX\[-5\] _06927_ rbzero.debug_overlay.playerX\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__o21ai_1
XFILLER_184_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11486_ rbzero.tex_g1\[3\] _03729_ _03730_ _03652_ vssd1 vssd1 vccd1 vccd1 _04269_
+ sky130_fd_sc_hd__a31o_1
XFILLER_183_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16013_ _08617_ _08626_ vssd1 vssd1 vccd1 vccd1 _08627_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_0__02751_ _02751_ vssd1 vssd1 vccd1 vccd1 clknet_0__02751_ sky130_fd_sc_hd__clkbuf_16
X_13225_ _05945_ _05944_ _05981_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__and3_1
X_10437_ rbzero.tex_b0\[49\] rbzero.tex_b0\[48\] _03280_ vssd1 vssd1 vccd1 vccd1 _03284_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13156_ _05491_ _05616_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__nand2_1
X_10368_ rbzero.tex_b1\[17\] rbzero.tex_b1\[18\] _03243_ vssd1 vssd1 vccd1 vccd1 _03248_
+ sky130_fd_sc_hd__mux2_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _04849_ _04867_ _04868_ _04843_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__o211a_1
XFILLER_151_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13087_ _05827_ _05828_ _05839_ _05843_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__o2bb2a_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17964_ _02182_ vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10299_ rbzero.tex_b1\[50\] rbzero.tex_b1\[51\] _03210_ vssd1 vssd1 vccd1 vccd1 _03212_
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19703_ clknet_leaf_74_i_clk _00634_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12038_ _03524_ _03461_ _03459_ _03469_ _04790_ net35 vssd1 vssd1 vccd1 vccd1 _04811_
+ sky130_fd_sc_hd__mux4_1
X_16915_ rbzero.wall_tracer.trackDistX\[7\] rbzero.wall_tracer.stepDistX\[7\] vssd1
+ vssd1 vccd1 vccd1 _09522_ sky130_fd_sc_hd__nand2_1
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17895_ _02146_ vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19634_ clknet_leaf_59_i_clk _00565_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16846_ _09444_ _09451_ vssd1 vssd1 vccd1 vccd1 _09453_ sky130_fd_sc_hd__nor2_1
X_19145__308 clknet_1_1__leaf__02746_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__inv_2
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19565_ clknet_leaf_36_i_clk _00496_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16777_ _09376_ _09384_ vssd1 vssd1 vccd1 vccd1 _09385_ sky130_fd_sc_hd__xnor2_1
X_13989_ _06734_ vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__clkbuf_1
X_18516_ _02475_ vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15728_ _08388_ _08410_ vssd1 vssd1 vccd1 vccd1 _08411_ sky130_fd_sc_hd__xnor2_1
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19496_ clknet_leaf_47_i_clk _00442_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[3\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_179_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15659_ _08206_ _08341_ vssd1 vssd1 vccd1 vccd1 _08342_ sky130_fd_sc_hd__xnor2_1
XFILLER_178_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18378_ rbzero.pov.spi_counter\[6\] rbzero.pov.spi_counter\[5\] _02426_ vssd1 vssd1
+ vccd1 vccd1 _02431_ sky130_fd_sc_hd__nand3_1
XFILLER_159_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17329_ _01651_ _09709_ rbzero.wall_tracer.trackDistY\[9\] _01523_ vssd1 vssd1 vccd1
+ vccd1 _00580_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_146_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19039__213 clknet_1_0__leaf__02735_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__inv_2
XFILLER_147_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20340_ net400 _01271_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20271_ net331 _01202_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__02740_ clknet_0__02740_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02740_
+ sky130_fd_sc_hd__clkbuf_16
X_19011__187 clknet_1_1__leaf__02733_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__inv_2
XFILLER_84_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19085__255 clknet_1_1__leaf__02739_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__inv_2
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_75 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_75/HI o_rgb[2] sky130_fd_sc_hd__conb_1
XFILLER_71_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_86 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_86/HI o_rgb[17] sky130_fd_sc_hd__conb_1
X_11340_ _04076_ _04091_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__nor2_1
Xtop_ew_algofoogle_97 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_97/HI zeros[6] sky130_fd_sc_hd__conb_1
XFILLER_193_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11271_ _03782_ _04051_ _04055_ _04040_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__and4bb_4
X_20469_ net125 _01400_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[60\] sky130_fd_sc_hd__dfxtp_1
X_13010_ _05732_ _05757_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__xnor2_1
X_10222_ _03171_ vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10153_ rbzero.tex_g0\[56\] rbzero.tex_g0\[55\] _03132_ vssd1 vssd1 vccd1 vccd1 _03135_
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10084_ rbzero.tex_g1\[24\] rbzero.tex_g1\[25\] _03095_ vssd1 vssd1 vccd1 vccd1 _03099_
+ sky130_fd_sc_hd__mux2_1
X_14961_ _07628_ _07627_ vssd1 vssd1 vccd1 vccd1 _07649_ sky130_fd_sc_hd__and2b_1
XFILLER_121_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16700_ rbzero.wall_tracer.trackDistX\[5\] rbzero.wall_tracer.stepDistX\[5\] vssd1
+ vssd1 vccd1 vccd1 _09309_ sky130_fd_sc_hd__nor2_1
XFILLER_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13912_ _06664_ _06665_ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__nand2_1
X_17680_ _01942_ _01945_ _01953_ vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__o21ai_1
X_14892_ _07533_ _07577_ _07578_ _07579_ vssd1 vssd1 vccd1 vccd1 _07580_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16631_ _09227_ _09239_ vssd1 vssd1 vccd1 vccd1 _09240_ sky130_fd_sc_hd__xnor2_1
X_13843_ _06593_ _06599_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__xnor2_2
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19350_ _02828_ _02829_ _02830_ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__a21o_1
X_16562_ _09164_ _09171_ vssd1 vssd1 vccd1 vccd1 _09172_ sky130_fd_sc_hd__xnor2_2
XFILLER_16_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13774_ _06517_ _06523_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10986_ _03770_ _03771_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__nand2_1
XFILLER_16_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18301_ rbzero.spi_registers.spi_buffer\[4\] rbzero.spi_registers.new_leak\[4\] _02379_
+ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__mux2_1
X_15513_ _08195_ _08196_ vssd1 vssd1 vccd1 vccd1 _08197_ sky130_fd_sc_hd__nor2_1
X_12725_ _05465_ _05479_ _05450_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__or3b_1
X_19281_ _02767_ _02768_ _02769_ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__o21ai_1
XFILLER_71_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16493_ _08643_ _07960_ _08071_ _08107_ vssd1 vssd1 vccd1 vccd1 _09103_ sky130_fd_sc_hd__o22a_1
XFILLER_128_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18232_ _03338_ _02342_ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__or2_1
X_15444_ _08024_ _08023_ vssd1 vssd1 vccd1 vccd1 _08129_ sky130_fd_sc_hd__or2b_1
XFILLER_188_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12656_ _05409_ _05410_ _05411_ _05412_ _05333_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__a221oi_1
XFILLER_90_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18163_ rbzero.map_overlay.i_mapdy\[0\] _02292_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__or2_1
X_11607_ _04315_ _04388_ _03830_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__mux2_1
X_12587_ _05158_ _05253_ _05311_ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__mux2_1
X_15375_ rbzero.wall_tracer.texu\[2\] _06853_ _08059_ _08060_ _03498_ vssd1 vssd1
+ vccd1 vccd1 _00477_ sky130_fd_sc_hd__o221a_1
XFILLER_168_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17114_ _09529_ _09702_ _09700_ vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__a21oi_2
X_14326_ _07011_ _07012_ _07013_ vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__o21ai_2
XFILLER_183_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11538_ rbzero.tex_b0\[63\] _04155_ _04156_ _03611_ vssd1 vssd1 vccd1 vccd1 _04320_
+ sky130_fd_sc_hd__a31o_1
X_18094_ net42 rbzero.spi_registers.ss_buffer\[0\] _03337_ vssd1 vssd1 vccd1 vccd1
+ _02252_ sky130_fd_sc_hd__mux2_1
XFILLER_143_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17045_ _09636_ _09649_ vssd1 vssd1 vccd1 vccd1 _09650_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11469_ rbzero.tex_g1\[27\] _03729_ _03730_ _03652_ vssd1 vssd1 vccd1 vccd1 _04252_
+ sky130_fd_sc_hd__a31o_1
X_14257_ rbzero.wall_tracer.visualWallDist\[-5\] _06944_ rbzero.wall_tracer.state\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__mux2_1
XFILLER_87_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__02734_ _02734_ vssd1 vssd1 vccd1 vccd1 clknet_0__02734_ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13208_ _05880_ _05928_ _05964_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__or3_1
XFILLER_87_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14188_ _06858_ _06866_ _06873_ _06875_ vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__or4_4
XFILLER_125_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13139_ _05895_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__inv_2
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17947_ _02173_ vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__clkbuf_1
XFILLER_97_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17878_ _02122_ _02133_ _02134_ _02123_ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__a31o_1
X_16829_ _07993_ _08333_ vssd1 vssd1 vccd1 vccd1 _09436_ sky130_fd_sc_hd__nor2_1
XFILLER_26_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19617_ clknet_leaf_39_i_clk _00548_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19548_ clknet_leaf_37_i_clk _00479_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19479_ clknet_leaf_49_i_clk _00425_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20323_ net383 _01254_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20254_ net314 _01185_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20185_ net245 _01116_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09996_ _03052_ vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_90_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02723_ clknet_0__02723_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__02723_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_56_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10840_ rbzero.row_render.texu\[2\] rbzero.row_render.texu\[1\] _03624_ _03625_ vssd1
+ vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__or4_1
XFILLER_44_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10771_ _03546_ _03549_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12510_ _05246_ _05251_ _05266_ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__and3_1
X_13490_ _06001_ _05995_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__nor2_1
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12441_ _05193_ _05197_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__or2_1
XFILLER_200_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18913__99 clknet_1_1__leaf__02723_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__inv_2
X_15160_ _07724_ _07833_ _07846_ vssd1 vssd1 vccd1 vccd1 _07847_ sky130_fd_sc_hd__a21oi_1
X_12372_ rbzero.wall_tracer.visualWallDist\[-5\] _05067_ _03487_ vssd1 vssd1 vccd1
+ vccd1 _05129_ sky130_fd_sc_hd__a21o_1
XFILLER_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_126_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18996__175 clknet_1_1__leaf__02730_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__inv_2
X_11323_ rbzero.debug_overlay.vplaneY\[-3\] _04092_ _04090_ rbzero.debug_overlay.vplaneY\[-8\]
+ _04107_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__a221o_1
X_14111_ rbzero.wall_tracer.stepDistX\[-7\] _06679_ _00008_ vssd1 vssd1 vccd1 vccd1
+ _06820_ sky130_fd_sc_hd__mux2_1
XFILLER_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15091_ _07776_ _07777_ vssd1 vssd1 vccd1 vccd1 _07779_ sky130_fd_sc_hd__and2_1
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11254_ _03503_ _04038_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__or2_1
X_14042_ _05210_ _05334_ _06736_ _06774_ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__o31ai_4
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10205_ _03162_ vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18850_ rbzero.pov.ready_buffer\[6\] _02635_ _02687_ _02672_ vssd1 vssd1 vccd1 vccd1
+ _01065_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_58_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_192_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11185_ rbzero.tex_r1\[13\] _03919_ _03768_ _03673_ vssd1 vssd1 vccd1 vccd1 _03970_
+ sky130_fd_sc_hd__a31o_1
XFILLER_133_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17801_ _02062_ _02063_ _02064_ _02065_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__a211o_1
X_10136_ net48 rbzero.tex_g0\[63\] _03050_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__mux2_1
XFILLER_121_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18781_ rbzero.debug_overlay.facingX\[-1\] _02645_ vssd1 vssd1 vccd1 vccd1 _02650_
+ sky130_fd_sc_hd__and2_1
XFILLER_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15993_ _07265_ _08191_ vssd1 vssd1 vccd1 vccd1 _08607_ sky130_fd_sc_hd__nor2_1
XFILLER_67_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17732_ _02001_ rbzero.wall_tracer.rayAddendX\[2\] vssd1 vssd1 vccd1 vccd1 _02002_
+ sky130_fd_sc_hd__xnor2_1
X_14944_ _07616_ _07631_ _07619_ vssd1 vssd1 vccd1 vccd1 _07632_ sky130_fd_sc_hd__o21a_1
X_10067_ rbzero.tex_g1\[32\] rbzero.tex_g1\[33\] _03084_ vssd1 vssd1 vccd1 vccd1 _03090_
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17663_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.debug_overlay.vplaneX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__or2_1
X_14875_ _07550_ _07561_ _07562_ vssd1 vssd1 vccd1 vccd1 _07563_ sky130_fd_sc_hd__a21oi_1
XFILLER_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19402_ rbzero.traced_texVinit\[8\] _02868_ _08454_ _08716_ vssd1 vssd1 vccd1 vccd1
+ _01436_ sky130_fd_sc_hd__a22o_1
X_16614_ _07984_ _08316_ vssd1 vssd1 vccd1 vccd1 _09223_ sky130_fd_sc_hd__nand2_1
X_13826_ _06581_ _06582_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__nor2_1
XFILLER_90_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17594_ _01879_ vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__clkbuf_1
X_19333_ _02812_ _02814_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__nand2_1
XFILLER_188_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16545_ _09046_ _09050_ vssd1 vssd1 vccd1 vccd1 _09155_ sky130_fd_sc_hd__or2_1
XFILLER_62_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13757_ _06485_ _06494_ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10969_ rbzero.tex_r0\[53\] rbzero.tex_r0\[52\] _03690_ vssd1 vssd1 vccd1 vccd1 _03755_
+ sky130_fd_sc_hd__mux2_1
X_12708_ _05356_ _05459_ _05460_ _05464_ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__a31o_2
X_19264_ rbzero.traced_texa\[-11\] rbzero.texV\[-11\] vssd1 vssd1 vccd1 vccd1 _02761_
+ sky130_fd_sc_hd__or2_1
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16476_ _09082_ _09083_ _09084_ vssd1 vssd1 vccd1 vccd1 _09087_ sky130_fd_sc_hd__a21o_1
XFILLER_148_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13688_ _06392_ _06444_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__or2b_1
XFILLER_188_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18215_ _03338_ _02330_ vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__or2_1
X_15427_ _08110_ _08111_ vssd1 vssd1 vccd1 vccd1 _08112_ sky130_fd_sc_hd__nor2_1
XFILLER_176_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12639_ _05238_ _05242_ _05311_ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__mux2_1
XFILLER_129_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18146_ _03901_ _02287_ _02258_ _03852_ vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__and4b_2
XFILLER_156_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15358_ _08042_ _08043_ vssd1 vssd1 vccd1 vccd1 _08044_ sky130_fd_sc_hd__nor2_2
XFILLER_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14309_ _06993_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__buf_4
XFILLER_171_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18077_ _02242_ vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15289_ _07853_ _07973_ _07974_ vssd1 vssd1 vccd1 vccd1 _07975_ sky130_fd_sc_hd__a21o_1
XFILLER_172_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17028_ _09281_ _09534_ vssd1 vssd1 vccd1 vccd1 _09633_ sky130_fd_sc_hd__nor2_1
XFILLER_176_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09850_ rbzero.tex_r1\[5\] rbzero.tex_r1\[6\] _02965_ vssd1 vssd1 vccd1 vccd1 _02974_
+ sky130_fd_sc_hd__mux2_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09781_ rbzero.tex_r1\[38\] rbzero.tex_r1\[39\] _02932_ vssd1 vssd1 vccd1 vccd1 _02938_
+ sky130_fd_sc_hd__mux2_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19123__288 clknet_1_0__leaf__02744_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__inv_2
XFILLER_33_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19197__356 clknet_1_0__leaf__02750_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__inv_2
XFILLER_167_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20306_ net366 _01237_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20237_ net297 _01168_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19017__193 clknet_1_0__leaf__02733_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__inv_2
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20168_ net228 _01099_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09979_ _03043_ vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _05516_ _05593_ _05728_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__or3_1
X_20099_ clknet_leaf_88_i_clk _01030_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ _03911_ _04666_ _04685_ _04686_ net42 vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__a32o_1
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _07346_ _07347_ vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__nor2_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _03524_ _03461_ _03838_ _02901_ net9 net10 vssd1 vssd1 vccd1 vccd1 _04648_
+ sky130_fd_sc_hd__mux4_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _06121_ _05991_ vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__nor2_1
X_10823_ _03558_ _03603_ _03608_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__or3b_1
X_14591_ _07274_ _07276_ _07277_ vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__a21oi_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16330_ _08940_ _08941_ vssd1 vssd1 vccd1 vccd1 _08942_ sky130_fd_sc_hd__nor2_1
XFILLER_38_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13542_ _06245_ _06298_ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__nor2_1
XFILLER_197_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10754_ _03539_ rbzero.row_render.wall\[1\] vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__nor2_1
XFILLER_111_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16261_ _08871_ _08872_ vssd1 vssd1 vccd1 vccd1 _08873_ sky130_fd_sc_hd__nor2_1
XFILLER_13_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13473_ _05902_ vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__buf_2
X_10685_ rbzero.wall_tracer.state\[11\] vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__inv_2
XFILLER_71_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18000_ _02201_ vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__clkbuf_1
X_15212_ _07185_ _07757_ _07898_ vssd1 vssd1 vccd1 vccd1 _07899_ sky130_fd_sc_hd__nor3_1
XFILLER_139_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12424_ _05153_ _05163_ _05177_ _05179_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__o211ai_2
XFILLER_199_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16192_ _07213_ _08682_ vssd1 vssd1 vccd1 vccd1 _08805_ sky130_fd_sc_hd__or2_2
XFILLER_139_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15143_ _07803_ _07804_ vssd1 vssd1 vccd1 vccd1 _07830_ sky130_fd_sc_hd__or2b_2
X_12355_ rbzero.debug_overlay.facingX\[-9\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__or2_1
XFILLER_142_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11306_ _03463_ _04040_ _04062_ _04052_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__or4_2
X_19951_ net180 _00882_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[31\] sky130_fd_sc_hd__dfxtp_1
X_15074_ _07185_ _07748_ _07756_ _07199_ _07761_ vssd1 vssd1 vccd1 vccd1 _07762_ sky130_fd_sc_hd__o41a_1
X_12286_ rbzero.debug_overlay.facingX\[-7\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__nand2_1
XFILLER_141_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11237_ _03840_ _03520_ _03834_ _04021_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__and4_1
X_18902_ _02722_ vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__clkbuf_1
X_14025_ rbzero.wall_tracer.stepDistY\[5\] _06765_ _06718_ vssd1 vssd1 vccd1 vccd1
+ _06766_ sky130_fd_sc_hd__mux2_1
X_19882_ clknet_leaf_23_i_clk _00813_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_136_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11168_ rbzero.tex_r1\[35\] _03733_ _03952_ _03666_ vssd1 vssd1 vccd1 vccd1 _03953_
+ sky130_fd_sc_hd__o211a_1
XFILLER_121_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18833_ _02081_ _02635_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__nand2_1
XFILLER_68_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10119_ _03072_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__buf_4
Xclkbuf_0__02433_ _02433_ vssd1 vssd1 vccd1 vccd1 clknet_0__02433_ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18764_ rbzero.debug_overlay.facingX\[-8\] _02638_ vssd1 vssd1 vccd1 vccd1 _02640_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11099_ _03879_ _03880_ _03883_ _03884_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__a211o_1
X_15976_ _08562_ _08589_ _08590_ _08522_ vssd1 vssd1 vccd1 vccd1 _08591_ sky130_fd_sc_hd__a31o_1
XFILLER_110_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17715_ _01985_ rbzero.wall_tracer.rayAddendX\[1\] vssd1 vssd1 vccd1 vccd1 _01986_
+ sky130_fd_sc_hd__nand2_1
X_14927_ _07594_ _07596_ vssd1 vssd1 vccd1 vccd1 _07615_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18695_ _02582_ _02584_ _02585_ _02586_ vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__o211a_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17646_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.wall_tracer.rayAddendX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__or2_1
X_14858_ _07410_ _07543_ vssd1 vssd1 vccd1 vccd1 _07546_ sky130_fd_sc_hd__and2_1
XFILLER_91_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13809_ _06561_ _06564_ _06565_ vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__a21o_1
X_17577_ _01847_ _01850_ _01848_ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__a21boi_1
XFILLER_63_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14789_ _07475_ _07476_ vssd1 vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__nor2b_2
XFILLER_95_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19316_ _02800_ _02801_ _02802_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__a21o_1
XFILLER_189_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16528_ _09136_ _09137_ vssd1 vssd1 vccd1 vccd1 _09138_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16459_ _09068_ _09069_ vssd1 vssd1 vccd1 vccd1 _09070_ sky130_fd_sc_hd__nor2_1
XFILLER_164_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18129_ _04828_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__buf_2
XFILLER_191_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09902_ rbzero.tex_r0\[47\] rbzero.tex_r0\[46\] _02995_ vssd1 vssd1 vccd1 vccd1 _03003_
+ sky130_fd_sc_hd__mux2_1
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20022_ clknet_leaf_88_i_clk _00953_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09833_ _02909_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__clkbuf_4
XFILLER_58_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09764_ rbzero.tex_r1\[46\] rbzero.tex_r1\[47\] _02921_ vssd1 vssd1 vccd1 vccd1 _02929_
+ sky130_fd_sc_hd__mux2_1
XFILLER_100_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18431__71 clknet_1_0__leaf__02438_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__inv_2
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19205__363 clknet_1_1__leaf__02751_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__inv_2
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10470_ rbzero.tex_b0\[33\] rbzero.tex_b0\[32\] _03291_ vssd1 vssd1 vccd1 vccd1 _03301_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12140_ _04890_ _04897_ _04898_ _04901_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__or4bb_1
XFILLER_151_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12071_ _04836_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__buf_4
XFILLER_150_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11022_ _03772_ _03807_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__nand2_1
XFILLER_110_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15830_ rbzero.traced_texa\[9\] _08463_ _08462_ rbzero.wall_tracer.visualWallDist\[9\]
+ vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__a22o_1
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _03526_ _03501_ vssd1 vssd1 vccd1 vccd1 _08441_ sky130_fd_sc_hd__or2_1
X_12973_ _05516_ _05728_ _05593_ _05729_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__or4b_1
XFILLER_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ _01781_ _01780_ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__and2b_1
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14712_ _07377_ _07379_ _07378_ _06901_ vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__a22o_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18480_ rbzero.pov.spi_buffer\[10\] rbzero.pov.spi_buffer\[11\] _02455_ vssd1 vssd1
+ vccd1 vccd1 _02457_ sky130_fd_sc_hd__mux2_1
X_11924_ net25 net26 _04690_ _04698_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__o31a_2
X_15692_ _08373_ _08374_ vssd1 vssd1 vccd1 vccd1 _08375_ sky130_fd_sc_hd__nand2_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.wall_tracer.rayAddendY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__or2_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _07254_ _07258_ _07253_ vssd1 vssd1 vccd1 vccd1 _07331_ sky130_fd_sc_hd__a21bo_1
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ net42 _04622_ _04623_ _04630_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__a31o_1
XFILLER_45_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10806_ rbzero.texV\[5\] _03561_ _03559_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__a21oi_2
X_17362_ _01673_ vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14574_ _07251_ _07252_ _07261_ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__o21ai_2
X_11786_ net19 vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__inv_2
XFILLER_198_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16313_ _08799_ _08924_ vssd1 vssd1 vccd1 vccd1 _08925_ sky130_fd_sc_hd__xor2_1
X_13525_ _06192_ _06210_ vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__nor2_1
XFILLER_159_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10737_ gpout0.hpos\[3\] vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__clkbuf_4
X_17293_ _08512_ _01620_ _01527_ vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__a21o_1
XFILLER_201_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19032_ clknet_1_1__leaf__02732_ vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__buf_1
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16244_ _08854_ _08855_ vssd1 vssd1 vccd1 vccd1 _08856_ sky130_fd_sc_hd__nor2_1
XFILLER_186_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13456_ _05768_ _06098_ _06106_ vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__a21oi_1
X_10668_ gpout0.hpos\[4\] vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__inv_2
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ rbzero.wall_tracer.visualWallDist\[8\] vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__inv_2
X_16175_ _08672_ _08674_ _08673_ vssd1 vssd1 vccd1 vccd1 _08788_ sky130_fd_sc_hd__a21bo_1
X_13387_ _06037_ _06036_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__xnor2_1
X_10599_ rbzero.map_rom.f4 vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__clkbuf_4
XFILLER_126_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15126_ rbzero.debug_overlay.playerY\[-7\] rbzero.debug_overlay.playerX\[-7\] _06850_
+ vssd1 vssd1 vccd1 vccd1 _07814_ sky130_fd_sc_hd__mux2_1
XFILLER_126_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12338_ _05037_ _05046_ _05035_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__a21bo_1
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19934_ net163 _00865_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[14\] sky130_fd_sc_hd__dfxtp_1
X_15057_ _07100_ _07138_ vssd1 vssd1 vccd1 vccd1 _07745_ sky130_fd_sc_hd__nor2_1
X_12269_ _04929_ _05025_ vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__nand2_1
XFILLER_96_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14008_ _05315_ _06750_ _05376_ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__a21o_1
X_19865_ clknet_leaf_24_i_clk _00796_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_95_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18816_ rbzero.pov.ready_buffer\[12\] _02663_ _02669_ _02643_ vssd1 vssd1 vccd1 vccd1
+ _01049_ sky130_fd_sc_hd__o211a_1
XFILLER_56_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19796_ clknet_leaf_18_i_clk _00727_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_49_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18747_ rbzero.debug_overlay.playerY\[4\] _02619_ _02411_ vssd1 vssd1 vccd1 vccd1
+ _02626_ sky130_fd_sc_hd__o21ai_1
X_15959_ _08485_ _08573_ _08574_ _08507_ _08575_ vssd1 vssd1 vccd1 vccd1 _08576_ sky130_fd_sc_hd__o311a_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18678_ rbzero.pov.ready_buffer\[71\] _02540_ _02571_ _02572_ _02543_ vssd1 vssd1
+ vccd1 vccd1 _02573_ sky130_fd_sc_hd__o221a_1
XFILLER_93_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17629_ _04932_ _04942_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__or2_1
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20005_ clknet_leaf_91_i_clk _00936_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_09816_ _02956_ vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09747_ rbzero.tex_r1\[54\] rbzero.tex_r1\[55\] _02910_ vssd1 vssd1 vccd1 vccd1 _02920_
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19129__294 clknet_1_1__leaf__02744_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__inv_2
XFILLER_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ rbzero.tex_b1\[58\] _03663_ _03823_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__a21o_1
XFILLER_30_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11571_ rbzero.tex_b0\[22\] _03617_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__and2_1
XFILLER_23_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13310_ _06038_ _06065_ _06066_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__a21oi_1
XFILLER_195_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10522_ _03328_ vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14290_ _06977_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__clkbuf_4
XFILLER_155_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10453_ _03292_ vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__clkbuf_1
X_13241_ _05989_ _05993_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__xnor2_1
XFILLER_196_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10384_ _03256_ vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__clkbuf_1
X_13172_ _05880_ _05928_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__nor2_1
XFILLER_151_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12123_ _04877_ _04878_ _04883_ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__or3b_1
XFILLER_112_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17980_ rbzero.pov.spi_buffer\[43\] rbzero.pov.ready_buffer\[43\] _02186_ vssd1 vssd1
+ vccd1 vccd1 _02191_ sky130_fd_sc_hd__mux2_1
XFILLER_46_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16931_ _09490_ _09491_ _09493_ vssd1 vssd1 vccd1 vccd1 _09537_ sky130_fd_sc_hd__o21ai_2
X_12054_ net34 _04779_ net35 _04780_ _04826_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__o41a_2
XFILLER_117_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11005_ _03788_ _03789_ _03790_ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__a21oi_1
X_16862_ _09269_ _09467_ vssd1 vssd1 vccd1 vccd1 _09469_ sky130_fd_sc_hd__or2_1
X_19650_ clknet_leaf_45_i_clk _00581_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15813_ _08447_ vssd1 vssd1 vccd1 vccd1 _08460_ sky130_fd_sc_hd__clkbuf_4
X_18601_ rbzero.pov.spi_buffer\[68\] rbzero.pov.spi_buffer\[69\] _02510_ vssd1 vssd1
+ vccd1 vccd1 _02520_ sky130_fd_sc_hd__mux2_1
X_19581_ clknet_leaf_62_i_clk _00512_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
X_16793_ _09210_ _09297_ _09295_ vssd1 vssd1 vccd1 vccd1 _09401_ sky130_fd_sc_hd__a21o_1
XFILLER_77_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18532_ rbzero.pov.spi_buffer\[35\] rbzero.pov.spi_buffer\[36\] _02477_ vssd1 vssd1
+ vccd1 vccd1 _02484_ sky130_fd_sc_hd__mux2_1
XFILLER_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15744_ _08424_ _08426_ vssd1 vssd1 vccd1 vccd1 _08427_ sky130_fd_sc_hd__nor2_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12956_ _05701_ _05712_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__xnor2_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ rbzero.pov.spi_buffer\[2\] rbzero.pov.spi_buffer\[3\] _02444_ vssd1 vssd1
+ vccd1 vccd1 _02448_ sky130_fd_sc_hd__mux2_1
XFILLER_34_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11907_ net24 _04670_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__and2b_1
X_15675_ _08244_ _08254_ _08256_ vssd1 vssd1 vccd1 vccd1 _08358_ sky130_fd_sc_hd__a21bo_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _05630_ _05643_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__xnor2_1
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _01702_ _01712_ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__xnor2_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18410__52 clknet_1_1__leaf__02436_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__inv_2
X_14626_ _07312_ _07313_ vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__nand2_1
XFILLER_60_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _04612_ net62 _04613_ net13 vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__o211a_1
XFILLER_61_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ rbzero.spi_registers.new_mapd\[1\] rbzero.spi_registers.spi_buffer\[1\] _01663_
+ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__mux2_1
X_14557_ _07209_ _07243_ vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__and2_1
XFILLER_60_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11769_ net7 _04510_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__nand2_1
XFILLER_140_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13508_ _06260_ _06263_ vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__nor2_1
X_17276_ _01602_ _01603_ _01604_ vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__and3_1
XFILLER_158_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14488_ _07175_ _04949_ _03492_ _07171_ vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__or4_2
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16227_ _08836_ _08837_ _08592_ _08596_ vssd1 vssd1 vccd1 vccd1 _08840_ sky130_fd_sc_hd__a211o_1
X_13439_ _05616_ _05768_ _06056_ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__and3_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16158_ _07993_ _07857_ vssd1 vssd1 vccd1 vccd1 _08771_ sky130_fd_sc_hd__nor2_1
XFILLER_138_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15109_ _07287_ _07781_ _07795_ vssd1 vssd1 vccd1 vccd1 _07797_ sky130_fd_sc_hd__and3_1
XFILLER_177_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16089_ _08355_ _08419_ _08417_ vssd1 vssd1 vccd1 vccd1 _08703_ sky130_fd_sc_hd__a21o_1
XFILLER_170_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19917_ clknet_leaf_95_i_clk _00848_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19848_ clknet_leaf_24_i_clk _00779_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_110_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19779_ clknet_leaf_83_i_clk _00710_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20485_ clknet_leaf_38_i_clk _01416_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12810_ _05556_ _05566_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__xnor2_1
X_13790_ _06439_ _06545_ _05557_ _05904_ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__o211ai_1
XFILLER_76_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _05492_ _05497_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__xor2_1
XFILLER_43_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19062__234 clknet_1_0__leaf__02737_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__inv_2
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _04950_ _08141_ _06860_ _06787_ vssd1 vssd1 vccd1 vccd1 _08145_ sky130_fd_sc_hd__and4bb_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12672_ _05270_ _05427_ _05428_ _05356_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__o31a_1
XFILLER_179_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__04486_ clknet_0__04486_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04486_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _07096_ _07098_ vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__xnor2_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11623_ rbzero.tex_b1\[47\] rbzero.tex_b1\[46\] _04188_ vssd1 vssd1 vccd1 vccd1 _04404_
+ sky130_fd_sc_hd__mux2_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15391_ _07853_ _07973_ vssd1 vssd1 vccd1 vccd1 _08076_ sky130_fd_sc_hd__nand2_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17130_ _01461_ _01473_ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__xnor2_2
XFILLER_156_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14342_ _04928_ _07028_ _07029_ vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__a21oi_1
XFILLER_196_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11554_ rbzero.tex_b0\[38\] _03617_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__and2_1
XFILLER_195_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17061_ _09664_ _09665_ vssd1 vssd1 vccd1 vccd1 _09666_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10505_ _03319_ vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14273_ rbzero.debug_overlay.playerX\[-4\] rbzero.debug_overlay.playerX\[-5\] _06927_
+ vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__or3_1
X_11485_ rbzero.tex_g1\[2\] _03664_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__and2_1
XFILLER_155_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16012_ _08624_ _08625_ vssd1 vssd1 vccd1 vccd1 _08626_ sky130_fd_sc_hd__nor2_1
XFILLER_13_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__02750_ _02750_ vssd1 vssd1 vccd1 vccd1 clknet_0__02750_ sky130_fd_sc_hd__clkbuf_16
X_13224_ _05942_ _05980_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__xor2_1
XFILLER_100_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10436_ _03283_ vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13155_ _05606_ _05861_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__nand2_1
XFILLER_98_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10367_ _03247_ vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__clkbuf_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _04846_ _04844_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__or2b_1
X_10298_ _03211_ vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__clkbuf_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17963_ rbzero.pov.spi_buffer\[35\] rbzero.pov.ready_buffer\[35\] _02175_ vssd1 vssd1
+ vccd1 vccd1 _02182_ sky130_fd_sc_hd__mux2_1
X_13086_ _05823_ _05842_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__nor2_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19702_ clknet_leaf_73_i_clk _00633_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12037_ _04792_ _04807_ _04808_ _04809_ _04798_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__a221o_1
X_16914_ rbzero.wall_tracer.trackDistX\[7\] rbzero.wall_tracer.stepDistX\[7\] vssd1
+ vssd1 vccd1 vccd1 _09521_ sky130_fd_sc_hd__nor2_1
X_17894_ rbzero.pov.spi_buffer\[2\] rbzero.pov.ready_buffer\[2\] _02143_ vssd1 vssd1
+ vccd1 vccd1 _02146_ sky130_fd_sc_hd__mux2_1
XFILLER_93_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19633_ clknet_leaf_53_i_clk _00564_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16845_ _09444_ _09451_ vssd1 vssd1 vccd1 vccd1 _09452_ sky130_fd_sc_hd__and2_1
XFILLER_66_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16776_ _09269_ _09383_ vssd1 vssd1 vccd1 vccd1 _09384_ sky130_fd_sc_hd__xnor2_1
X_19564_ clknet_leaf_63_i_clk _00495_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13988_ rbzero.wall_tracer.stepDistY\[0\] _06733_ _06718_ vssd1 vssd1 vccd1 vccd1
+ _06734_ sky130_fd_sc_hd__mux2_1
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15727_ _08407_ _08409_ vssd1 vssd1 vccd1 vccd1 _08410_ sky130_fd_sc_hd__xor2_2
X_18515_ rbzero.pov.spi_buffer\[27\] rbzero.pov.spi_buffer\[28\] _02466_ vssd1 vssd1
+ vccd1 vccd1 _02475_ sky130_fd_sc_hd__mux2_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12939_ _05517_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__inv_2
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19495_ clknet_leaf_47_i_clk _00441_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_33_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15658_ _07084_ _07270_ _08339_ _08340_ vssd1 vssd1 vccd1 vccd1 _08341_ sky130_fd_sc_hd__o31a_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14609_ _07117_ _07156_ _07215_ _07296_ _07214_ vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__o32a_1
X_18377_ rbzero.pov.spi_counter\[5\] _02426_ rbzero.pov.spi_counter\[6\] vssd1 vssd1
+ vccd1 vccd1 _02430_ sky130_fd_sc_hd__a21o_1
XFILLER_57_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15589_ _08265_ _08272_ vssd1 vssd1 vccd1 vccd1 _08273_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17328_ _01649_ _01650_ _01522_ vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__o21a_1
XFILLER_105_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17259_ rbzero.wall_tracer.trackDistY\[0\] rbzero.wall_tracer.stepDistY\[0\] vssd1
+ vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__or2_1
XFILLER_146_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20270_ net330 _01201_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_76 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_76/HI o_rgb[3] sky130_fd_sc_hd__conb_1
XFILLER_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_87 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_87/HI o_rgb[18] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_98 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_98/HI zeros[7] sky130_fd_sc_hd__conb_1
XFILLER_192_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20468_ net148 _01399_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[59\] sky130_fd_sc_hd__dfxtp_1
X_11270_ _04052_ _04054_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__nor2_1
XFILLER_106_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10221_ rbzero.tex_g0\[24\] rbzero.tex_g0\[23\] _03166_ vssd1 vssd1 vccd1 vccd1 _03171_
+ sky130_fd_sc_hd__mux2_1
X_20399_ net459 _01330_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10152_ _03134_ vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10083_ _03098_ vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__clkbuf_1
X_14960_ _06873_ _07617_ _07647_ vssd1 vssd1 vccd1 vccd1 _07648_ sky130_fd_sc_hd__or3_1
XFILLER_48_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13911_ _05324_ _06609_ _06644_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__a21o_1
XFILLER_102_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14891_ _06872_ _06933_ vssd1 vssd1 vccd1 vccd1 _07579_ sky130_fd_sc_hd__or2_1
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16630_ _09237_ _09238_ vssd1 vssd1 vccd1 vccd1 _09239_ sky130_fd_sc_hd__nor2_1
XFILLER_47_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13842_ _06575_ _06586_ _06584_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__a21oi_1
XFILLER_56_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16561_ _09169_ _09170_ vssd1 vssd1 vccd1 vccd1 _09171_ sky130_fd_sc_hd__nor2_1
XFILLER_62_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13773_ _06504_ _06512_ _06529_ vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__a21oi_1
XFILLER_62_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18927__112 clknet_1_1__leaf__02724_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__inv_2
X_10985_ rbzero.row_render.size\[1\] rbzero.row_render.size\[0\] vssd1 vssd1 vccd1
+ vccd1 _03771_ sky130_fd_sc_hd__nor2_1
XFILLER_90_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15512_ _07265_ _07960_ _08070_ _07269_ vssd1 vssd1 vccd1 vccd1 _08196_ sky130_fd_sc_hd__o22a_1
XFILLER_71_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18300_ _02383_ vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__clkbuf_1
X_12724_ _05477_ _05480_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__nand2_1
X_19280_ _02772_ _02773_ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__nand2_1
X_16492_ _09101_ vssd1 vssd1 vccd1 vccd1 _09102_ sky130_fd_sc_hd__inv_2
XFILLER_167_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18231_ rbzero.color_floor\[3\] rbzero.spi_registers.new_floor\[3\] _02335_ vssd1
+ vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__mux2_1
X_15443_ _08116_ _08127_ vssd1 vssd1 vccd1 vccd1 _08128_ sky130_fd_sc_hd__xor2_1
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12655_ _05261_ _05349_ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__nand2_1
XFILLER_169_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11606_ _03764_ _04349_ _04384_ _04387_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__a31o_1
XFILLER_50_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18162_ rbzero.spi_registers.new_mapd\[15\] _02290_ _02298_ _02275_ vssd1 vssd1 vccd1
+ vccd1 _00766_ sky130_fd_sc_hd__o211a_1
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15374_ _07937_ _08057_ _08058_ _04832_ vssd1 vssd1 vccd1 vccd1 _08060_ sky130_fd_sc_hd__a31o_1
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12586_ _05339_ _05342_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__or2_1
X_17113_ _09615_ _09619_ _09706_ _09716_ vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__a31o_1
X_14325_ _06856_ _06872_ vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__or2_1
XFILLER_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11537_ rbzero.tex_b0\[62\] _03617_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__and2_1
X_18093_ _02251_ vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17044_ _09641_ _09648_ vssd1 vssd1 vccd1 vccd1 _09649_ sky130_fd_sc_hd__xnor2_1
XFILLER_144_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14256_ rbzero.debug_overlay.playerY\[-5\] _06943_ _04927_ vssd1 vssd1 vccd1 vccd1
+ _06944_ sky130_fd_sc_hd__mux2_1
X_11468_ rbzero.tex_g1\[26\] _03664_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__and2_1
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__02733_ _02733_ vssd1 vssd1 vccd1 vccd1 clknet_0__02733_ sky130_fd_sc_hd__clkbuf_16
X_13207_ _05928_ _05963_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__nor2_1
X_10419_ _03274_ vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__clkbuf_1
X_14187_ _06874_ vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__buf_2
XFILLER_139_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11399_ _04181_ _04182_ _03635_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__mux2_1
XFILLER_87_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18973__154 clknet_1_0__leaf__02728_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__inv_2
XFILLER_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _05646_ _05686_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__nor2_1
XFILLER_112_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13069_ _05697_ _05480_ _05820_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__and3_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17946_ rbzero.pov.spi_buffer\[27\] rbzero.pov.ready_buffer\[27\] _02164_ vssd1 vssd1
+ vccd1 vccd1 _02173_ sky130_fd_sc_hd__mux2_1
XFILLER_100_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17877_ rbzero.spi_registers.spi_counter\[4\] _02129_ vssd1 vssd1 vccd1 vccd1 _02134_
+ sky130_fd_sc_hd__or2_1
XFILLER_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19616_ clknet_leaf_60_i_clk _00547_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16828_ _09325_ _09433_ _09434_ vssd1 vssd1 vccd1 vccd1 _09435_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19547_ clknet_leaf_30_i_clk _00478_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16759_ _09021_ _09256_ _09255_ _09253_ vssd1 vssd1 vccd1 vccd1 _09367_ sky130_fd_sc_hd__o31a_1
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19478_ clknet_leaf_49_i_clk _00424_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20322_ net382 _01253_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20253_ net313 _01184_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19091__260 clknet_1_0__leaf__02740_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__inv_2
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20184_ net244 _01115_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09995_ rbzero.tex_r0\[3\] rbzero.tex_r0\[2\] _03050_ vssd1 vssd1 vccd1 vccd1 _03052_
+ sky130_fd_sc_hd__mux2_1
XFILLER_142_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18438__77 clknet_1_1__leaf__02439_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__inv_2
XFILLER_131_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10770_ _03552_ _03555_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__or2_2
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12440_ _05194_ _05196_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__xnor2_2
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12371_ _05037_ _05046_ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__xnor2_2
XFILLER_201_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19174__335 clknet_1_1__leaf__02748_ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__inv_2
XFILLER_181_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14110_ _06819_ vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_138_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11322_ rbzero.debug_overlay.vplaneY\[-4\] _04089_ _04085_ rbzero.debug_overlay.vplaneY\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__a22o_1
X_15090_ _07776_ _07777_ vssd1 vssd1 vccd1 vccd1 _07778_ sky130_fd_sc_hd__nor2_1
XFILLER_180_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14041_ _06778_ vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__clkbuf_1
X_11253_ gpout0.hpos\[3\] _04033_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__nor2_1
XFILLER_140_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10204_ rbzero.tex_g0\[32\] rbzero.tex_g0\[31\] _03155_ vssd1 vssd1 vccd1 vccd1 _03162_
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11184_ rbzero.tex_r1\[15\] _03664_ _03968_ _03677_ vssd1 vssd1 vccd1 vccd1 _03969_
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17800_ rbzero.wall_tracer.rayAddendX\[6\] rbzero.wall_tracer.rayAddendX\[5\] rbzero.wall_tracer.rayAddendX\[4\]
+ rbzero.wall_tracer.rayAddendX\[3\] _02000_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__o41a_1
X_10135_ _03125_ vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__clkbuf_1
X_15992_ _08376_ _08357_ vssd1 vssd1 vccd1 vccd1 _08606_ sky130_fd_sc_hd__or2b_1
X_18780_ rbzero.pov.ready_buffer\[40\] _02636_ _02649_ _02643_ vssd1 vssd1 vccd1 vccd1
+ _01033_ sky130_fd_sc_hd__o211a_1
XFILLER_0_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14943_ _07620_ vssd1 vssd1 vccd1 vccd1 _07631_ sky130_fd_sc_hd__inv_2
X_10066_ _03089_ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__clkbuf_1
X_17731_ _02000_ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__clkbuf_4
XFILLER_134_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14874_ _07560_ _07551_ vssd1 vssd1 vccd1 vccd1 _07562_ sky130_fd_sc_hd__and2b_1
X_17662_ _01936_ _01937_ _03485_ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__o21ai_1
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19401_ rbzero.traced_texVinit\[7\] _02868_ _08431_ _01745_ vssd1 vssd1 vccd1 vccd1
+ _01435_ sky130_fd_sc_hd__a22o_1
XFILLER_75_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16613_ _09220_ _09221_ vssd1 vssd1 vccd1 vccd1 _09222_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13825_ _06222_ _06580_ vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__and2_1
XFILLER_169_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17593_ rbzero.wall_tracer.rayAddendY\[8\] _01878_ _03509_ vssd1 vssd1 vccd1 vccd1
+ _01879_ sky130_fd_sc_hd__mux2_1
XFILLER_51_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16544_ _09037_ _09040_ _09034_ vssd1 vssd1 vccd1 vccd1 _09154_ sky130_fd_sc_hd__a21bo_1
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19332_ rbzero.traced_texa\[1\] rbzero.texV\[1\] vssd1 vssd1 vccd1 vccd1 _02817_
+ sky130_fd_sc_hd__nand2_1
X_13756_ _05862_ _06230_ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__nor2_1
X_10968_ _03674_ _03749_ _03753_ _03679_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__a211o_1
XFILLER_188_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12707_ _05367_ _05350_ _05462_ _05323_ _05463_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__a221o_1
XFILLER_149_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19263_ rbzero.traced_texa\[-11\] rbzero.texV\[-11\] vssd1 vssd1 vccd1 vccd1 _02760_
+ sky130_fd_sc_hd__nand2_1
X_16475_ _09085_ vssd1 vssd1 vccd1 vccd1 _09086_ sky130_fd_sc_hd__inv_2
XFILLER_188_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13687_ _06346_ _06391_ vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__or2_1
X_10899_ _03684_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__buf_6
X_15426_ _08106_ _08109_ vssd1 vssd1 vccd1 vccd1 _08111_ sky130_fd_sc_hd__and2_1
X_18214_ rbzero.color_sky\[4\] rbzero.spi_registers.new_sky\[4\] _02320_ vssd1 vssd1
+ vccd1 vccd1 _02330_ sky130_fd_sc_hd__mux2_1
X_12638_ _05274_ _05329_ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__nor2_4
XFILLER_157_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15357_ _08040_ _08041_ vssd1 vssd1 vccd1 vccd1 _08043_ sky130_fd_sc_hd__and2_1
X_18145_ gpout0.vpos\[2\] gpout0.vpos\[1\] _02286_ vssd1 vssd1 vccd1 vccd1 _02287_
+ sky130_fd_sc_hd__and3_1
XFILLER_200_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12569_ _05256_ _05228_ _05231_ _05219_ _05324_ _05325_ vssd1 vssd1 vccd1 vccd1 _05326_
+ sky130_fd_sc_hd__mux4_1
XFILLER_157_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14308_ _06941_ _06995_ vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__xnor2_1
X_18076_ rbzero.spi_registers.spi_buffer\[14\] rbzero.spi_registers.spi_buffer\[13\]
+ _02226_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__mux2_1
X_15288_ _06856_ _07084_ _07235_ _06874_ vssd1 vssd1 vccd1 vccd1 _07974_ sky130_fd_sc_hd__o22a_1
XFILLER_172_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17027_ _09532_ _09535_ _09631_ vssd1 vssd1 vccd1 vccd1 _09632_ sky130_fd_sc_hd__a21o_1
X_14239_ rbzero.debug_overlay.playerX\[-6\] _06888_ vssd1 vssd1 vccd1 vccd1 _06927_
+ sky130_fd_sc_hd__or2_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _02937_ vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__clkbuf_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17929_ _02142_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__buf_4
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20305_ net365 _01236_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20236_ net296 _01167_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20167_ net227 _01098_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[14\] sky130_fd_sc_hd__dfxtp_1
X_09978_ rbzero.tex_r0\[11\] rbzero.tex_r0\[10\] _03039_ vssd1 vssd1 vccd1 vccd1 _03043_
+ sky130_fd_sc_hd__mux2_1
XFILLER_104_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20098_ clknet_leaf_90_i_clk _01029_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-6\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11940_ _04670_ _04714_ net24 vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__and3b_1
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ net12 net11 _04646_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__and3_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _06121_ _05987_ _06366_ vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__nor3_1
X_10822_ _03556_ _03557_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__nand2_1
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14590_ _07274_ _07276_ _07277_ vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__and3_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13541_ _06001_ _06071_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__nor2_1
X_10753_ rbzero.row_render.wall\[0\] vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__clkinv_2
XFILLER_186_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16260_ _08864_ _08870_ vssd1 vssd1 vccd1 vccd1 _08872_ sky130_fd_sc_hd__nor2_1
XFILLER_200_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13472_ _06183_ _06185_ vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__xnor2_1
XFILLER_186_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10684_ _02904_ _03468_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__nand2_2
XFILLER_139_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15211_ _07178_ _07897_ vssd1 vssd1 vccd1 vccd1 _07898_ sky130_fd_sc_hd__or2_1
XFILLER_127_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12423_ _05159_ _05176_ _05163_ _05179_ _05153_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__a311o_1
XFILLER_200_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16191_ _07213_ _07185_ _07199_ _08803_ vssd1 vssd1 vccd1 vccd1 _08804_ sky130_fd_sc_hd__a31o_1
XFILLER_127_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15142_ rbzero.wall_tracer.texu\[0\] _06853_ _07828_ _07829_ _03498_ vssd1 vssd1
+ vccd1 vccd1 _00475_ sky130_fd_sc_hd__o221a_1
X_12354_ rbzero.wall_tracer.visualWallDist\[-9\] _05066_ rbzero.wall_tracer.rcp_sel\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__a21o_1
XFILLER_181_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11305_ _04073_ _04080_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__nor2_4
X_19950_ net179 _00881_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[30\] sky130_fd_sc_hd__dfxtp_1
X_15073_ _07155_ _07180_ vssd1 vssd1 vccd1 vccd1 _07761_ sky130_fd_sc_hd__or2b_1
X_12285_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__nand2_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14024_ _06630_ _06764_ vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__or2_1
X_18901_ _02707_ _02721_ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__and2_1
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11236_ gpout0.vpos\[5\] _03517_ _04020_ _03524_ vssd1 vssd1 vccd1 vccd1 _04021_
+ sky130_fd_sc_hd__nor4_1
X_19881_ clknet_leaf_22_i_clk _00812_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18832_ rbzero.pov.ready_buffer\[19\] _02663_ _02678_ _02672_ vssd1 vssd1 vccd1 vccd1
+ _01056_ sky130_fd_sc_hd__o211a_1
X_11167_ rbzero.tex_r1\[34\] _03767_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__or2_1
X_10118_ _03116_ vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__clkbuf_1
X_18417__58 clknet_1_1__leaf__02437_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__inv_2
X_18763_ rbzero.pov.ready_buffer\[33\] _02636_ _02639_ _02586_ vssd1 vssd1 vccd1 vccd1
+ _01026_ sky130_fd_sc_hd__o211a_1
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11098_ gpout0.vpos\[5\] rbzero.map_overlay.i_othery\[2\] vssd1 vssd1 vccd1 vccd1
+ _03884_ sky130_fd_sc_hd__xor2_1
X_15975_ _08586_ _08587_ _08588_ vssd1 vssd1 vccd1 vccd1 _08590_ sky130_fd_sc_hd__o21ai_1
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17714_ rbzero.debug_overlay.vplaneX\[10\] vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__buf_2
X_14926_ _07601_ _07603_ vssd1 vssd1 vccd1 vccd1 _07614_ sky130_fd_sc_hd__xnor2_1
X_10049_ _03080_ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18694_ _04828_ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__clkbuf_4
XFILLER_64_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17645_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.wall_tracer.rayAddendX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__nand2_1
XFILLER_64_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14857_ _07517_ _07519_ vssd1 vssd1 vccd1 vccd1 _07545_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13808_ _06331_ _06432_ _06335_ vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__and3_1
XFILLER_90_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17576_ _01861_ _01862_ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__nand2_1
X_14788_ _07472_ _07474_ vssd1 vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__nand2_1
XFILLER_189_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19315_ _02800_ _02801_ _02802_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__nand3_1
XFILLER_177_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16527_ _08899_ _07857_ vssd1 vssd1 vccd1 vccd1 _09137_ sky130_fd_sc_hd__nor2_1
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13739_ _06461_ _06479_ _06495_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__and3_1
XFILLER_17_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16458_ _09066_ _09067_ vssd1 vssd1 vccd1 vccd1 _09069_ sky130_fd_sc_hd__and2_1
XFILLER_31_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15409_ _07983_ _07985_ _07987_ vssd1 vssd1 vccd1 vccd1 _08094_ sky130_fd_sc_hd__o21ai_1
XFILLER_129_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16389_ _08998_ _08999_ vssd1 vssd1 vccd1 vccd1 _09000_ sky130_fd_sc_hd__nor2_1
XFILLER_145_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18128_ rbzero.map_overlay.i_othery\[2\] _02268_ vssd1 vssd1 vccd1 vccd1 _02274_
+ sky130_fd_sc_hd__or2_1
XFILLER_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18059_ _02233_ vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09901_ _03002_ vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20021_ clknet_leaf_94_i_clk _00952_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_98_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09832_ _02964_ vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09763_ _02928_ vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_86_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_42_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_57_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_167_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12070_ net72 rbzero.wall_tracer.state\[9\] _02907_ vssd1 vssd1 vccd1 vccd1 _04836_
+ sky130_fd_sc_hd__and3_2
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11021_ _03770_ _03771_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__or2_1
X_20219_ net279 _01150_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15760_ _08440_ vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__clkbuf_1
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _05495_ _05727_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__xor2_1
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ _07396_ _07398_ vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__nand2_1
X_11923_ net22 _04693_ _04695_ _04697_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__a31o_1
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15691_ _08364_ _08372_ vssd1 vssd1 vccd1 vccd1 _08374_ sky130_fd_sc_hd__or2_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _07325_ _07319_ vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__or2b_1
X_17430_ rbzero.debug_overlay.vplaneY\[-3\] rbzero.wall_tracer.rayAddendY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__and2_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ net12 _04624_ _04629_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__and3_1
XFILLER_60_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _03588_ _03590_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__nand2_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14573_ _07259_ _07260_ vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__nand2_1
X_17361_ rbzero.spi_registers.new_mapd\[9\] rbzero.spi_registers.spi_buffer\[9\] _01662_
+ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__mux2_1
XFILLER_198_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11785_ _04554_ _04557_ _04561_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__and3_1
XFILLER_198_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16312_ _07662_ _08803_ vssd1 vssd1 vccd1 vccd1 _08924_ sky130_fd_sc_hd__nor2_1
X_13524_ _06278_ _06280_ vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__nand2_1
XFILLER_14_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10736_ _03514_ _03516_ _03521_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__nor3_4
X_17292_ _01618_ _01619_ vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__xnor2_1
XFILLER_198_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16243_ _08730_ _08734_ _08732_ vssd1 vssd1 vccd1 vccd1 _08855_ sky130_fd_sc_hd__a21oi_1
X_13455_ _06056_ _06200_ _06197_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__and3_1
XFILLER_51_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10667_ gpout0.hpos\[3\] vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__inv_2
XFILLER_142_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12406_ _03488_ _05078_ _05162_ _05080_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__o31a_2
X_16174_ _08664_ _08666_ _08663_ vssd1 vssd1 vccd1 vccd1 _08787_ sky130_fd_sc_hd__a21bo_1
XFILLER_51_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13386_ _05862_ _06035_ vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__nor2_1
X_10598_ _03373_ _03352_ _03393_ _03343_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__a22o_1
X_15125_ _07700_ _07702_ vssd1 vssd1 vccd1 vccd1 _07813_ sky130_fd_sc_hd__xor2_4
X_12337_ _03488_ _05091_ _05092_ _05093_ vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_142_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19933_ net162 _00864_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[13\] sky130_fd_sc_hd__dfxtp_1
X_15056_ _07730_ _07742_ _07743_ vssd1 vssd1 vccd1 vccd1 _07744_ sky130_fd_sc_hd__o21ai_2
X_12268_ _04929_ _05025_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__or2_1
X_14007_ _06588_ _06598_ _06605_ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__a21o_1
X_11219_ _03915_ _04003_ _03830_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__mux2_1
XFILLER_122_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19864_ clknet_leaf_25_i_clk _00795_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12199_ rbzero.wall_tracer.trackDistY\[3\] vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__inv_2
XFILLER_95_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18815_ rbzero.debug_overlay.vplaneX\[-8\] _02660_ vssd1 vssd1 vccd1 vccd1 _02669_
+ sky130_fd_sc_hd__or2_1
XFILLER_110_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19795_ clknet_leaf_18_i_clk _00726_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18746_ _02582_ _02624_ rbzero.debug_overlay.playerY\[4\] vssd1 vssd1 vccd1 vccd1
+ _02625_ sky130_fd_sc_hd__o21a_1
X_15958_ _04946_ _08174_ vssd1 vssd1 vccd1 vccd1 _08575_ sky130_fd_sc_hd__nand2_1
XFILLER_110_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14909_ _07588_ _07593_ vssd1 vssd1 vccd1 vccd1 _07597_ sky130_fd_sc_hd__nor2_1
XFILLER_36_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18677_ rbzero.debug_overlay.playerX\[3\] _02566_ _02412_ vssd1 vssd1 vccd1 vccd1
+ _02572_ sky130_fd_sc_hd__a21o_1
X_15889_ rbzero.wall_tracer.trackDistX\[-11\] rbzero.wall_tracer.stepDistX\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _08514_ sky130_fd_sc_hd__or2_1
XFILLER_36_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17628_ _01907_ vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17559_ _01845_ _01846_ _01834_ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__a21o_1
XFILLER_149_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09815_ rbzero.tex_r1\[22\] rbzero.tex_r1\[23\] _02954_ vssd1 vssd1 vccd1 vccd1 _02956_
+ sky130_fd_sc_hd__mux2_1
X_20004_ clknet_leaf_91_i_clk _00935_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09746_ _02919_ vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11570_ _04350_ _04351_ _03740_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__mux2_1
XFILLER_156_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10521_ rbzero.tex_b0\[9\] rbzero.tex_b0\[8\] _03324_ vssd1 vssd1 vccd1 vccd1 _03328_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13240_ _05989_ _05993_ _05996_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__and3_1
XFILLER_196_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10452_ rbzero.tex_b0\[42\] rbzero.tex_b0\[41\] _03291_ vssd1 vssd1 vccd1 vccd1 _03292_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13171_ _05493_ _05517_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__or2_1
X_10383_ rbzero.tex_b1\[10\] rbzero.tex_b1\[11\] _03254_ vssd1 vssd1 vccd1 vccd1 _03256_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12122_ _04877_ _04878_ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__o21bai_1
XFILLER_123_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16930_ _09532_ _09535_ vssd1 vssd1 vccd1 vccd1 _09536_ sky130_fd_sc_hd__xnor2_1
X_12053_ _04782_ _04785_ _04789_ _04825_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__a31o_2
XFILLER_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11004_ rbzero.row_render.size\[6\] _03466_ _03777_ _02900_ vssd1 vssd1 vccd1 vccd1
+ _03790_ sky130_fd_sc_hd__o22ai_1
XFILLER_89_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16861_ _09269_ _09467_ vssd1 vssd1 vccd1 vccd1 _09468_ sky130_fd_sc_hd__nand2_1
XFILLER_42_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18600_ _02519_ vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__clkbuf_1
X_15812_ rbzero.traced_texa\[-5\] _08457_ _08459_ rbzero.wall_tracer.visualWallDist\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__a22o_1
X_19580_ clknet_leaf_66_i_clk _00511_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
X_16792_ _09320_ _09399_ vssd1 vssd1 vccd1 vccd1 _09400_ sky130_fd_sc_hd__xnor2_1
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18531_ _02483_ vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__clkbuf_1
X_15743_ _08289_ _08291_ _08425_ vssd1 vssd1 vccd1 vccd1 _08426_ sky130_fd_sc_hd__o21a_1
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12955_ _05709_ _05710_ _05711_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__o21ai_2
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11906_ net25 _04678_ _04679_ _04680_ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__a211o_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18462_ _02447_ vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15674_ _08228_ _08238_ _08236_ vssd1 vssd1 vccd1 vccd1 _08357_ sky130_fd_sc_hd__a21o_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ _05641_ _05642_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__nor2_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _01703_ _01710_ _01711_ vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__a21boi_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14625_ _07302_ _07310_ _07311_ vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__nand3_1
X_11837_ _04612_ _04314_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__nand2_1
X_18393_ clknet_1_1__leaf__02433_ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__buf_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14556_ _07209_ _07243_ vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__nor2_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _01664_ vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11768_ _04540_ _04541_ _04545_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__o21ai_1
XFILLER_186_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13507_ _06260_ _06263_ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__xor2_1
X_10719_ rbzero.wall_tracer.state\[14\] _03506_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__nand2_1
X_17275_ _01602_ _01603_ _01604_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__a21o_1
X_14487_ _06787_ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__inv_2
XFILLER_186_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11699_ rbzero.row_render.texu\[3\] rbzero.row_render.texu\[2\] _03539_ rbzero.row_render.side
+ _02899_ _03783_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__mux4_1
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13438_ _05480_ _06098_ _06106_ _06086_ vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__a211o_1
X_16226_ _08838_ vssd1 vssd1 vccd1 vccd1 _08839_ sky130_fd_sc_hd__inv_2
XFILLER_173_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16157_ _08766_ _08767_ _08768_ _08769_ vssd1 vssd1 vccd1 vccd1 _08770_ sky130_fd_sc_hd__a31o_1
XFILLER_154_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13369_ _06125_ _06099_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__xnor2_1
XFILLER_182_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15108_ _07287_ _07781_ _07795_ vssd1 vssd1 vccd1 vccd1 _07796_ sky130_fd_sc_hd__a21oi_2
XFILLER_181_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16088_ _08636_ _08701_ vssd1 vssd1 vccd1 vccd1 _08702_ sky130_fd_sc_hd__xor2_1
XFILLER_103_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15039_ _07704_ _07726_ vssd1 vssd1 vccd1 vccd1 _07727_ sky130_fd_sc_hd__xnor2_1
X_19916_ clknet_leaf_0_i_clk _00847_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19847_ clknet_leaf_24_i_clk _00778_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_110_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19778_ clknet_leaf_82_i_clk _00709_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18729_ rbzero.debug_overlay.playerY\[0\] _07026_ rbzero.debug_overlay.playerY\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__o21ai_1
XFILLER_114_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20484_ clknet_leaf_38_i_clk _01415_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09729_ rbzero.tex_r1\[63\] net47 _02910_ vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__mux2_1
XFILLER_62_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12740_ _05493_ _05496_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__nor2_1
XFILLER_16_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _05329_ _05336_ _05337_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__and3_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _07097_ _06993_ vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__nor2_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11622_ rbzero.tex_b1\[45\] rbzero.tex_b1\[44\] _04189_ vssd1 vssd1 vccd1 vccd1 _04403_
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15390_ _07945_ _07947_ _07944_ vssd1 vssd1 vccd1 vccd1 _08075_ sky130_fd_sc_hd__a21bo_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ rbzero.debug_overlay.playerY\[-1\] _04928_ vssd1 vssd1 vccd1 vccd1 _07029_
+ sky130_fd_sc_hd__nor2_1
X_11553_ _03740_ _04332_ _04333_ _04334_ _03702_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__o221a_1
XFILLER_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17060_ _08862_ _08333_ vssd1 vssd1 vccd1 vccd1 _09665_ sky130_fd_sc_hd__nor2_1
X_10504_ rbzero.tex_b0\[17\] rbzero.tex_b0\[16\] _03313_ vssd1 vssd1 vccd1 vccd1 _03319_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14272_ rbzero.wall_tracer.visualWallDist\[-4\] _06959_ rbzero.wall_tracer.state\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__mux2_1
X_11484_ _04265_ _04266_ _03612_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__mux2_1
XFILLER_144_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16011_ _08618_ _08362_ _08623_ vssd1 vssd1 vccd1 vccd1 _08625_ sky130_fd_sc_hd__and3_1
XFILLER_137_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13223_ _05978_ _05979_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__nor2_1
X_10435_ rbzero.tex_b0\[50\] rbzero.tex_b0\[49\] _03280_ vssd1 vssd1 vccd1 vccd1 _03283_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13154_ _05875_ _05886_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__nand2_1
XFILLER_151_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10366_ rbzero.tex_b1\[18\] rbzero.tex_b1\[19\] _03243_ vssd1 vssd1 vccd1 vccd1 _03247_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12105_ _04853_ _04866_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__or2_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ _02181_ vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13085_ _05814_ _05816_ _05841_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__o21ai_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10297_ rbzero.tex_b1\[51\] rbzero.tex_b1\[52\] _03210_ vssd1 vssd1 vccd1 vccd1 _03211_
+ sky130_fd_sc_hd__mux2_1
X_19701_ clknet_leaf_74_i_clk _00632_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16913_ _09517_ _09518_ _09519_ vssd1 vssd1 vccd1 vccd1 _09520_ sky130_fd_sc_hd__o21ai_2
X_12036_ _04503_ _03902_ _04790_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__mux2_1
XFILLER_104_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17893_ _02145_ vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19632_ clknet_leaf_53_i_clk _00563_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
X_16844_ _09445_ _09450_ vssd1 vssd1 vccd1 vccd1 _09451_ sky130_fd_sc_hd__xor2_1
XFILLER_92_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19563_ clknet_leaf_36_i_clk _00494_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_16775_ _09379_ _09380_ _09382_ vssd1 vssd1 vccd1 vccd1 _09383_ sky130_fd_sc_hd__o21a_1
XFILLER_46_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13987_ _05390_ _06731_ _06732_ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__o21ai_4
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18514_ _02474_ vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__clkbuf_1
X_15726_ _08264_ _08275_ _08408_ vssd1 vssd1 vccd1 vccd1 _08409_ sky130_fd_sc_hd__a21oi_2
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ _05693_ _05694_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__and2b_1
X_19494_ clknet_leaf_52_i_clk _00440_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[1\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15657_ _08107_ _07257_ _07333_ _07084_ vssd1 vssd1 vccd1 vccd1 _08340_ sky130_fd_sc_hd__o22ai_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _05617_ _05625_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__xnor2_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14608_ rbzero.wall_tracer.visualWallDist\[-10\] _04839_ _06985_ _07114_ vssd1 vssd1
+ vccd1 vccd1 _07296_ sky130_fd_sc_hd__and4_1
X_18376_ rbzero.pov.spi_counter\[5\] _02426_ _02429_ vssd1 vssd1 vccd1 vccd1 _00849_
+ sky130_fd_sc_hd__o21a_1
X_15588_ _08145_ _08270_ _08271_ _08142_ vssd1 vssd1 vccd1 vccd1 _08272_ sky130_fd_sc_hd__a22oi_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17327_ _01646_ _01647_ _01648_ _03341_ vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__a31o_1
XFILLER_109_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14539_ _07218_ _07212_ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__or2b_1
XFILLER_146_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17258_ rbzero.wall_tracer.trackDistY\[0\] rbzero.wall_tracer.stepDistY\[0\] vssd1
+ vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__nand2_1
XFILLER_88_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16209_ _08636_ _08700_ _08699_ vssd1 vssd1 vccd1 vccd1 _08822_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17189_ _01524_ _01529_ _01530_ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__nand3b_1
XFILLER_143_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18950__133 clknet_1_1__leaf__02726_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__inv_2
XFILLER_111_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19046__219 clknet_1_1__leaf__02736_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__inv_2
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18386__30 clknet_1_0__leaf__02434_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__inv_2
XFILLER_25_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xtop_ew_algofoogle_77 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_77/HI o_rgb[4] sky130_fd_sc_hd__conb_1
XFILLER_137_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_88 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_88/HI o_rgb[19] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_99 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_99/HI zeros[8] sky130_fd_sc_hd__conb_1
XFILLER_123_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20467_ net147 _01398_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_180_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10220_ _03170_ vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20398_ net458 _01329_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[53\] sky130_fd_sc_hd__dfxtp_1
X_10151_ rbzero.tex_g0\[57\] rbzero.tex_g0\[56\] _03132_ vssd1 vssd1 vccd1 vccd1 _03134_
+ sky130_fd_sc_hd__mux2_1
XFILLER_121_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10082_ rbzero.tex_g1\[25\] rbzero.tex_g1\[26\] _03095_ vssd1 vssd1 vccd1 vccd1 _03098_
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13910_ _05380_ vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__clkbuf_4
X_14890_ _07101_ _07006_ _07048_ _07119_ vssd1 vssd1 vccd1 vccd1 _07578_ sky130_fd_sc_hd__o22a_1
XFILLER_130_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13841_ _06595_ _06597_ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__xor2_2
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16560_ _08805_ _09165_ _09168_ vssd1 vssd1 vccd1 vccd1 _09170_ sky130_fd_sc_hd__and3_1
X_13772_ _06337_ _06513_ _06528_ _06526_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__a31o_1
XFILLER_74_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10984_ rbzero.row_render.size\[2\] vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__inv_2
X_15511_ _08194_ vssd1 vssd1 vccd1 vccd1 _08195_ sky130_fd_sc_hd__inv_2
X_12723_ _05450_ _05479_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__xnor2_4
XFILLER_188_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16491_ _08643_ _08107_ _07960_ _08070_ vssd1 vssd1 vccd1 vccd1 _09101_ sky130_fd_sc_hd__or4_1
XFILLER_167_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18230_ _02341_ vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__clkbuf_1
X_15442_ _08125_ _08126_ vssd1 vssd1 vccd1 vccd1 _08127_ sky130_fd_sc_hd__and2_1
XFILLER_130_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12654_ _05242_ _05311_ _05338_ _05269_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__o211a_1
XFILLER_15_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11605_ _03642_ _04225_ _04386_ _03541_ _03537_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__o311a_1
XFILLER_168_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18161_ rbzero.map_overlay.i_mapdx\[5\] _02292_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__or2_1
XFILLER_184_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12585_ _05340_ _05341_ _05329_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__a21oi_1
X_15373_ _08057_ _08058_ _07937_ vssd1 vssd1 vccd1 vccd1 _08059_ sky130_fd_sc_hd__a21oi_1
X_17112_ _09613_ _09705_ _09704_ vssd1 vssd1 vccd1 vccd1 _09716_ sky130_fd_sc_hd__a21bo_1
X_14324_ _06875_ vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__clkbuf_4
X_11536_ _04316_ _04317_ _03740_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__mux2_1
XFILLER_129_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18092_ rbzero.spi_registers.mosi rbzero.spi_registers.mosi_buffer\[0\] _04834_ vssd1
+ vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__mux2_1
XFILLER_144_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17043_ _09646_ _09647_ vssd1 vssd1 vccd1 vccd1 _09648_ sky130_fd_sc_hd__nor2_1
X_14255_ _06942_ _06922_ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__xnor2_1
X_11467_ _04248_ _04249_ _03612_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__mux2_1
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__02732_ _02732_ vssd1 vssd1 vccd1 vccd1 clknet_0__02732_ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13206_ _05491_ _05962_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__nand2_1
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10418_ rbzero.tex_b0\[58\] rbzero.tex_b0\[57\] _03269_ vssd1 vssd1 vccd1 vccd1 _03274_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19151__314 clknet_1_0__leaf__02746_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__inv_2
X_14186_ rbzero.wall_tracer.visualWallDist\[2\] _06855_ vssd1 vssd1 vccd1 vccd1 _06874_
+ sky130_fd_sc_hd__nand2_2
X_11398_ rbzero.tex_g0\[11\] rbzero.tex_g0\[10\] _03662_ vssd1 vssd1 vccd1 vccd1 _04182_
+ sky130_fd_sc_hd__mux2_1
X_19239__14 clknet_1_0__leaf__02754_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__inv_2
XFILLER_180_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _05891_ _05893_ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__xnor2_1
X_10349_ rbzero.tex_b1\[26\] rbzero.tex_b1\[27\] _03232_ vssd1 vssd1 vccd1 vccd1 _03238_
+ sky130_fd_sc_hd__mux2_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _05802_ _05824_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__and2_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _02172_ vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__clkbuf_1
X_12019_ net34 vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__inv_2
XFILLER_79_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17876_ rbzero.spi_registers.spi_counter\[4\] _02129_ vssd1 vssd1 vccd1 vccd1 _02133_
+ sky130_fd_sc_hd__nand2_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19615_ clknet_leaf_61_i_clk _00546_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16827_ _08862_ _07961_ _08071_ _08888_ vssd1 vssd1 vccd1 vccd1 _09434_ sky130_fd_sc_hd__o22a_1
XFILLER_54_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19546_ clknet_leaf_41_i_clk _00477_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16758_ _09364_ _09365_ vssd1 vssd1 vccd1 vccd1 _09366_ sky130_fd_sc_hd__xor2_1
XFILLER_94_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15709_ _07646_ _08391_ vssd1 vssd1 vccd1 vccd1 _08392_ sky130_fd_sc_hd__or2_1
X_19477_ clknet_leaf_50_i_clk _00423_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16689_ _09210_ _09297_ vssd1 vssd1 vccd1 vccd1 _09298_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18359_ rbzero.pov.spi_counter\[1\] rbzero.pov.spi_counter\[0\] _02414_ vssd1 vssd1
+ vccd1 vccd1 _02417_ sky130_fd_sc_hd__and3_1
XFILLER_147_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20321_ net381 _01252_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20252_ net312 _01183_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09994_ _03051_ vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__clkbuf_1
X_20183_ net243 _01114_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12370_ _05120_ _05126_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__or2_1
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19100__268 clknet_1_0__leaf__02741_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__inv_2
XFILLER_193_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11321_ rbzero.debug_overlay.vplaneX\[10\] _04078_ _04105_ vssd1 vssd1 vccd1 vccd1
+ _04106_ sky130_fd_sc_hd__a21oi_2
X_20519_ clknet_leaf_24_i_clk _01450_ vssd1 vssd1 vccd1 vccd1 gpout1.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18957__139 clknet_1_0__leaf__02727_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__inv_2
XFILLER_180_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14040_ rbzero.wall_tracer.stepDistY\[8\] _06777_ _04836_ vssd1 vssd1 vccd1 vccd1
+ _06778_ sky130_fd_sc_hd__mux2_1
XFILLER_158_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11252_ _03513_ _04036_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__or2_1
X_10203_ _03161_ vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__clkbuf_1
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11183_ rbzero.tex_r1\[14\] _03620_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__or2_1
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10134_ rbzero.tex_g1\[0\] rbzero.tex_g1\[1\] _03117_ vssd1 vssd1 vccd1 vccd1 _03125_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15991_ _08375_ _08358_ vssd1 vssd1 vccd1 vccd1 _08605_ sky130_fd_sc_hd__or2b_1
XFILLER_47_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17730_ _01985_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__clkbuf_4
X_14942_ _07615_ _07629_ vssd1 vssd1 vccd1 vccd1 _07630_ sky130_fd_sc_hd__xor2_1
X_10065_ rbzero.tex_g1\[33\] rbzero.tex_g1\[34\] _03084_ vssd1 vssd1 vccd1 vccd1 _03089_
+ sky130_fd_sc_hd__mux2_1
XFILLER_134_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17661_ _01933_ _01934_ _01935_ vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__a21oi_1
X_14873_ _07551_ _07560_ vssd1 vssd1 vccd1 vccd1 _07561_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19400_ rbzero.traced_texVinit\[6\] _02868_ _08303_ _01745_ vssd1 vssd1 vccd1 vccd1
+ _01434_ sky130_fd_sc_hd__a22o_1
X_16612_ _09100_ _09104_ _09102_ vssd1 vssd1 vccd1 vccd1 _09221_ sky130_fd_sc_hd__a21oi_1
XFILLER_62_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13824_ _06222_ _06580_ vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__nor2_2
X_17592_ _01868_ _01869_ _01877_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__o21ai_1
XFILLER_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19331_ rbzero.traced_texa\[1\] rbzero.texV\[1\] vssd1 vssd1 vccd1 vccd1 _02816_
+ sky130_fd_sc_hd__or2_1
X_16543_ _09131_ _09152_ vssd1 vssd1 vccd1 vccd1 _09153_ sky130_fd_sc_hd__xnor2_2
XFILLER_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10967_ _03666_ _03750_ _03752_ _03670_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__o211a_1
X_13755_ _06497_ _06503_ _06502_ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__a21o_1
XFILLER_16_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12706_ _05325_ _05344_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__and2_1
X_19262_ _08439_ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__clkbuf_4
X_16474_ _09082_ _09083_ _09084_ vssd1 vssd1 vccd1 vccd1 _09085_ sky130_fd_sc_hd__and3_1
XFILLER_189_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10898_ _03603_ _03683_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__or2_4
X_13686_ _06440_ _06441_ _06442_ vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__nand3_1
XFILLER_188_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18213_ _02329_ vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__clkbuf_1
X_15425_ _08106_ _08109_ vssd1 vssd1 vccd1 vccd1 _08110_ sky130_fd_sc_hd__nor2_1
XFILLER_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12637_ _05367_ _05362_ _05393_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__a21o_1
XFILLER_19_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18144_ gpout0.vpos\[0\] _08450_ vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__and2_1
X_15356_ _08040_ _08041_ vssd1 vssd1 vccd1 vccd1 _08042_ sky130_fd_sc_hd__nor2_1
X_12568_ _05304_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__clkbuf_4
XFILLER_145_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11519_ rbzero.tex_g1\[47\] _03729_ _03730_ _03660_ vssd1 vssd1 vccd1 vccd1 _04302_
+ sky130_fd_sc_hd__a31o_1
X_14307_ _06972_ _06994_ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__xnor2_1
XFILLER_116_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18075_ _02241_ vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__clkbuf_1
X_15287_ _06874_ _07084_ vssd1 vssd1 vccd1 vccd1 _07973_ sky130_fd_sc_hd__nor2_1
XFILLER_8_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12499_ _05213_ _05214_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17026_ _09536_ _09560_ vssd1 vssd1 vccd1 vccd1 _09631_ sky130_fd_sc_hd__and2b_1
XFILLER_176_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14238_ rbzero.wall_tracer.visualWallDist\[-6\] _06925_ _03491_ vssd1 vssd1 vccd1
+ vccd1 _06926_ sky130_fd_sc_hd__mux2_1
XFILLER_109_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14169_ _06856_ vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__buf_2
XFILLER_124_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _02163_ vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__clkbuf_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17859_ rbzero.spi_registers.spi_counter\[2\] rbzero.spi_registers.spi_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__nor2_1
XFILLER_61_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19529_ clknet_leaf_66_i_clk _00001_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20304_ net364 _01235_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20235_ net295 _01166_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20166_ net226 _01097_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09977_ _03042_ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20097_ clknet_leaf_90_i_clk _01028_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_69_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ gpout0.hpos\[0\] _03527_ _03526_ _04020_ net9 net10 vssd1 vssd1 vccd1 vccd1
+ _04646_ sky130_fd_sc_hd__mux4_1
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19255__5 clknet_1_0__leaf__02433_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__inv_2
X_10821_ _03606_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__buf_6
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19180__340 clknet_1_1__leaf__02749_ vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__inv_2
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10752_ rbzero.row_render.side vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__inv_2
XFILLER_13_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13540_ _06008_ _06156_ vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__or2_1
XFILLER_158_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13471_ _06165_ _06190_ vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10683_ _03477_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__buf_6
XFILLER_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19024__199 clknet_1_1__leaf__02734_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__inv_2
X_12422_ _05080_ _05165_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__nand2_1
X_15210_ _04841_ rbzero.wall_tracer.stepDistX\[6\] _07895_ _07896_ vssd1 vssd1 vccd1
+ vccd1 _07897_ sky130_fd_sc_hd__o22ai_4
XFILLER_139_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16190_ _08681_ vssd1 vssd1 vccd1 vccd1 _08803_ sky130_fd_sc_hd__clkbuf_4
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12353_ _05067_ _04896_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__nor2_1
X_15141_ _07824_ _07827_ _04832_ vssd1 vssd1 vccd1 vccd1 _07829_ sky130_fd_sc_hd__a21o_1
XFILLER_126_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11304_ _04063_ _04070_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__nor2_4
X_15072_ _07749_ _07759_ vssd1 vssd1 vccd1 vccd1 _07760_ sky130_fd_sc_hd__xnor2_2
X_12284_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__nor2_1
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14023_ _06761_ _06762_ _06763_ _06711_ _05373_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__a32o_2
X_18900_ _03909_ _02719_ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__xnor2_1
X_11235_ _03523_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__clkbuf_4
X_19880_ clknet_leaf_23_i_clk _00811_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18831_ rbzero.debug_overlay.vplaneX\[-1\] _02660_ vssd1 vssd1 vccd1 vccd1 _02678_
+ sky130_fd_sc_hd__or2_1
XFILLER_84_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11166_ rbzero.tex_r1\[36\] _03919_ _03733_ _03950_ vssd1 vssd1 vccd1 vccd1 _03951_
+ sky130_fd_sc_hd__a31o_1
XFILLER_45_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10117_ rbzero.tex_g1\[8\] rbzero.tex_g1\[9\] _03106_ vssd1 vssd1 vccd1 vccd1 _03116_
+ sky130_fd_sc_hd__mux2_1
X_18762_ rbzero.debug_overlay.facingX\[-9\] _02638_ vssd1 vssd1 vccd1 vccd1 _02639_
+ sky130_fd_sc_hd__or2_1
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11097_ _03857_ rbzero.map_overlay.i_othery\[3\] _03881_ _03523_ _03882_ vssd1 vssd1
+ vccd1 vccd1 _03883_ sky130_fd_sc_hd__a221o_1
X_15974_ _08586_ _08587_ _08588_ vssd1 vssd1 vccd1 vccd1 _08589_ sky130_fd_sc_hd__or3_1
XFILLER_48_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17713_ _01984_ vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14925_ _07576_ _07605_ vssd1 vssd1 vccd1 vccd1 _07613_ sky130_fd_sc_hd__or2b_1
X_10048_ rbzero.tex_g1\[41\] rbzero.tex_g1\[42\] _03073_ vssd1 vssd1 vccd1 vccd1 _03080_
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18693_ _02583_ _02582_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__nand2_1
XFILLER_64_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17644_ rbzero.debug_overlay.vplaneX\[-9\] rbzero.wall_tracer.rayAddendX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__nand2_1
X_14856_ _07410_ _07543_ vssd1 vssd1 vccd1 vccd1 _07544_ sky130_fd_sc_hd__nor2_1
XFILLER_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13807_ _06332_ _06562_ _06563_ vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__a21o_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17575_ _01845_ _01859_ _01860_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__or3_1
XFILLER_95_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14787_ _07472_ _07474_ vssd1 vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__nor2_1
X_11999_ _04750_ _04393_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__nor2_1
XFILLER_16_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19314_ _02794_ _02797_ _02795_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__o21bai_1
X_16526_ _09134_ _09135_ vssd1 vssd1 vccd1 vccd1 _09136_ sky130_fd_sc_hd__nand2_1
XFILLER_91_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13738_ _06485_ _06494_ _06492_ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__a21o_1
XFILLER_56_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16457_ _09066_ _09067_ vssd1 vssd1 vccd1 vccd1 _09068_ sky130_fd_sc_hd__nor2_1
XFILLER_32_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13669_ _06382_ _06425_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__and2b_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15408_ _08066_ _08092_ vssd1 vssd1 vccd1 vccd1 _08093_ sky130_fd_sc_hd__xnor2_2
X_19176_ clknet_1_1__leaf__02743_ vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__buf_1
X_16388_ _08996_ _08997_ vssd1 vssd1 vccd1 vccd1 _08999_ sky130_fd_sc_hd__and2_1
XFILLER_157_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18127_ rbzero.spi_registers.new_other\[1\] _02264_ _02273_ _02266_ vssd1 vssd1 vccd1
+ vccd1 _00756_ sky130_fd_sc_hd__o211a_1
X_15339_ _08023_ _08024_ vssd1 vssd1 vccd1 vccd1 _08025_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18058_ rbzero.spi_registers.spi_buffer\[5\] rbzero.spi_registers.spi_buffer\[4\]
+ _02227_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__mux2_1
XFILLER_133_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17009_ _09613_ _09614_ vssd1 vssd1 vccd1 vccd1 _09615_ sky130_fd_sc_hd__nor2_2
X_09900_ rbzero.tex_r0\[48\] rbzero.tex_r0\[47\] _02995_ vssd1 vssd1 vccd1 vccd1 _03002_
+ sky130_fd_sc_hd__mux2_1
XFILLER_144_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20020_ clknet_leaf_94_i_clk _00951_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_09831_ rbzero.tex_r1\[14\] rbzero.tex_r1\[15\] _02954_ vssd1 vssd1 vccd1 vccd1 _02964_
+ sky130_fd_sc_hd__mux2_1
XFILLER_99_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09762_ rbzero.tex_r1\[47\] rbzero.tex_r1\[48\] _02921_ vssd1 vssd1 vccd1 vccd1 _02928_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11020_ _03773_ _03805_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__nand2_1
X_20218_ net278 _01149_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19212__369 clknet_1_0__leaf__02752_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__inv_2
XFILLER_77_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20149_ clknet_leaf_13_i_clk _01080_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _05697_ _05480_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__nand2_1
XFILLER_57_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14710_ _06998_ _07394_ _07397_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__o21ba_1
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ net22 _04696_ _04678_ net26 net25 vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__o2111ai_1
X_15690_ _08364_ _08372_ vssd1 vssd1 vccd1 vccd1 _08373_ sky130_fd_sc_hd__nand2_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _07291_ _07328_ vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__xor2_2
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ net49 _04622_ _04625_ net39 _04628_ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__a221o_1
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ _03586_ _03587_ rbzero.texV\[6\] vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__a21o_1
X_17360_ _01672_ vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__clkbuf_1
X_14572_ _07251_ _07252_ vssd1 vssd1 vccd1 vccd1 _07260_ sky130_fd_sc_hd__xor2_1
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11784_ net20 _04560_ net16 net17 vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__and4b_1
XFILLER_186_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16311_ _07877_ _08391_ vssd1 vssd1 vccd1 vccd1 _08923_ sky130_fd_sc_hd__or2_1
X_19106__274 clknet_1_1__leaf__02741_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__inv_2
XFILLER_185_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13523_ _06192_ _06279_ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__nor2_1
XFILLER_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10735_ _03517_ _03518_ _03519_ _03520_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__o31a_1
X_17291_ _01609_ _01613_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__nand2_1
XFILLER_186_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16242_ _08849_ _08853_ vssd1 vssd1 vccd1 vccd1 _08854_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13454_ _06192_ _06210_ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__and2_1
X_10666_ _03460_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__buf_2
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12405_ rbzero.wall_tracer.visualWallDist\[7\] _03480_ vssd1 vssd1 vccd1 vccd1 _05162_
+ sky130_fd_sc_hd__nor2_1
XFILLER_185_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16173_ _08764_ _08785_ vssd1 vssd1 vccd1 vccd1 _08786_ sky130_fd_sc_hd__xnor2_1
X_13385_ _06076_ _06141_ vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__or2_1
XFILLER_154_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10597_ _03391_ _03392_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__nand2_1
XFILLER_86_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15124_ _07810_ _07811_ vssd1 vssd1 vccd1 vccd1 _07812_ sky130_fd_sc_hd__nand2_1
XFILLER_127_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12336_ rbzero.wall_tracer.visualWallDist\[-3\] _05067_ _03487_ vssd1 vssd1 vccd1
+ vccd1 _05093_ sky130_fd_sc_hd__a21o_1
XFILLER_181_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19932_ net161 _00863_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15055_ _07119_ _07101_ _07136_ _07198_ vssd1 vssd1 vccd1 vccd1 _07743_ sky130_fd_sc_hd__or4_1
XFILLER_5_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12267_ rbzero.wall_tracer.mapY\[10\] _05024_ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11218_ _03537_ _03958_ _03995_ _04002_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__o31ai_2
X_14006_ _05376_ _06748_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__nand2_1
X_19863_ clknet_leaf_22_i_clk _00794_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12198_ rbzero.wall_tracer.trackDistY\[4\] vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__inv_2
XFILLER_150_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11149_ rbzero.tex_r1\[58\] _03926_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__or2_1
X_18814_ rbzero.pov.ready_buffer\[11\] _02666_ _02668_ _02651_ vssd1 vssd1 vccd1 vccd1
+ _01048_ sky130_fd_sc_hd__a211o_1
X_19794_ clknet_leaf_18_i_clk _00725_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18745_ _02607_ _02620_ vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__nor2_1
XFILLER_110_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15957_ _08570_ _08571_ _08572_ vssd1 vssd1 vccd1 vccd1 _08574_ sky130_fd_sc_hd__o21a_1
XFILLER_36_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14908_ _07579_ _07595_ vssd1 vssd1 vccd1 vccd1 _07596_ sky130_fd_sc_hd__xor2_1
XFILLER_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18676_ _02570_ vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__inv_2
XFILLER_64_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15888_ rbzero.wall_tracer.trackDistX\[-11\] rbzero.wall_tracer.stepDistX\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _08513_ sky130_fd_sc_hd__nand2_1
XFILLER_91_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17627_ _01906_ rbzero.map_rom.a6 _05009_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__mux2_1
XFILLER_63_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14839_ _07471_ _07526_ vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__nor2_1
XFILLER_36_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17558_ _01785_ _04109_ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__nand2_1
XFILLER_177_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16509_ _09112_ _09117_ vssd1 vssd1 vccd1 vccd1 _09119_ sky130_fd_sc_hd__nor2_1
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17489_ _01780_ _01781_ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20003_ clknet_leaf_92_i_clk _00934_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_09814_ _02955_ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09745_ rbzero.tex_r1\[55\] rbzero.tex_r1\[56\] _02910_ vssd1 vssd1 vccd1 vccd1 _02919_
+ sky130_fd_sc_hd__mux2_1
XFILLER_189_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10520_ _03327_ vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10451_ _03143_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__clkbuf_4
XFILLER_182_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13170_ _05484_ _05479_ _05472_ _05926_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__or4_2
XFILLER_108_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10382_ _03255_ vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12121_ _04880_ _04882_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__nand2_1
XFILLER_163_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12052_ net38 _04806_ _04819_ _04824_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__a31o_2
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11003_ rbzero.row_render.size\[6\] _03466_ _03781_ rbzero.row_render.size\[5\] vssd1
+ vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_78_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16860_ _09379_ _09466_ _09381_ vssd1 vssd1 vccd1 vccd1 _09467_ sky130_fd_sc_hd__o21a_1
XFILLER_131_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15811_ rbzero.traced_texa\[-6\] _08457_ _08459_ rbzero.wall_tracer.visualWallDist\[-6\]
+ vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__a22o_1
XFILLER_77_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16791_ _09396_ _09398_ vssd1 vssd1 vccd1 vccd1 _09399_ sky130_fd_sc_hd__xor2_1
XFILLER_120_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18530_ rbzero.pov.spi_buffer\[34\] rbzero.pov.spi_buffer\[35\] _02477_ vssd1 vssd1
+ vccd1 vccd1 _02483_ sky130_fd_sc_hd__mux2_1
X_15742_ _08292_ _08187_ vssd1 vssd1 vccd1 vccd1 _08425_ sky130_fd_sc_hd__or2b_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _05703_ _05708_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__or2b_1
XFILLER_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ rbzero.pov.spi_buffer\[1\] rbzero.pov.spi_buffer\[2\] _02444_ vssd1 vssd1
+ vccd1 vccd1 _02447_ sky130_fd_sc_hd__mux2_1
X_11905_ net26 vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__inv_2
X_15673_ _08281_ _08282_ vssd1 vssd1 vccd1 vccd1 _08356_ sky130_fd_sc_hd__or2_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _05631_ _05640_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__and2_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17412_ rbzero.debug_overlay.vplaneY\[-6\] rbzero.wall_tracer.rayAddendY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__nand2_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _07302_ _07310_ _07311_ vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__a21o_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ net9 vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__buf_2
XFILLER_61_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17343_ rbzero.spi_registers.new_mapd\[0\] rbzero.spi_registers.spi_buffer\[0\] _01663_
+ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__mux2_1
X_14555_ _07231_ _07242_ _07229_ vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _04496_ _04544_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__nand2_1
XFILLER_159_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13506_ _06173_ _06261_ _06262_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__a21boi_1
X_10718_ _03467_ _03503_ _03504_ _03505_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__and4b_4
X_17274_ _01595_ _01599_ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__nand2_1
XFILLER_146_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14486_ rbzero.wall_tracer.visualWallDist\[-10\] _06855_ vssd1 vssd1 vccd1 vccd1
+ _07174_ sky130_fd_sc_hd__and2_2
X_11698_ rbzero.row_render.texu\[1\] rbzero.row_render.texu\[0\] _02899_ vssd1 vssd1
+ vccd1 vccd1 _04478_ sky130_fd_sc_hd__mux2_1
X_16225_ _08592_ _08596_ _08836_ _08837_ vssd1 vssd1 vccd1 vccd1 _08838_ sky130_fd_sc_hd__o211a_1
XFILLER_139_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13437_ _06085_ _06094_ _06193_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__o21ai_1
X_10649_ _03433_ _03434_ _03435_ _03444_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__a211o_1
XFILLER_177_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16156_ _06858_ _07878_ _08000_ _07012_ vssd1 vssd1 vccd1 vccd1 _08769_ sky130_fd_sc_hd__o22a_1
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13368_ _05549_ _06055_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_41_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_15107_ _07793_ _07794_ vssd1 vssd1 vccd1 vccd1 _07795_ sky130_fd_sc_hd__nand2_1
XFILLER_170_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12319_ _05072_ _05075_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__nor2_1
X_16087_ _08699_ _08700_ vssd1 vssd1 vccd1 vccd1 _08701_ sky130_fd_sc_hd__and2b_1
XFILLER_138_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13299_ _06055_ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__buf_2
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15038_ _07724_ _07725_ vssd1 vssd1 vccd1 vccd1 _07726_ sky130_fd_sc_hd__nand2_1
X_19915_ clknet_leaf_0_i_clk _00846_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_111_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19846_ clknet_leaf_25_i_clk _00777_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16989_ _09496_ _09565_ _09594_ vssd1 vssd1 vccd1 vccd1 _09595_ sky130_fd_sc_hd__a21oi_1
XFILLER_3_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19777_ clknet_leaf_82_i_clk _00708_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18728_ rbzero.debug_overlay.playerY\[1\] rbzero.debug_overlay.playerY\[0\] _07026_
+ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__or3_1
XFILLER_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18659_ rbzero.pov.ready_buffer\[67\] _02411_ _02413_ _02557_ _02543_ vssd1 vssd1
+ vccd1 vccd1 _02558_ sky130_fd_sc_hd__o221a_1
XFILLER_184_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20483_ clknet_leaf_38_i_clk _01414_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_7_0_i_clk clknet_2_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_156_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09728_ _02909_ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__clkbuf_4
XFILLER_132_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _05338_ _05340_ _05341_ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__and3_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _04192_ _04399_ _04401_ _03702_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__o211a_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14340_ _07026_ _07027_ vssd1 vssd1 vccd1 vccd1 _07028_ sky130_fd_sc_hd__nand2_1
X_11552_ rbzero.tex_b0\[34\] _04247_ _03652_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__a21o_1
XFILLER_168_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10503_ _03318_ vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11483_ rbzero.tex_g1\[5\] rbzero.tex_g1\[4\] _04247_ vssd1 vssd1 vccd1 vccd1 _04266_
+ sky130_fd_sc_hd__mux2_1
X_14271_ rbzero.debug_overlay.playerY\[-4\] _06958_ _04927_ vssd1 vssd1 vccd1 vccd1
+ _06959_ sky130_fd_sc_hd__mux2_1
XFILLER_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16010_ _08618_ _08362_ _08623_ vssd1 vssd1 vccd1 vccd1 _08624_ sky130_fd_sc_hd__a21oi_1
XFILLER_100_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10434_ _03282_ vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13222_ _05936_ _05939_ _05977_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__and3_1
XFILLER_152_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19218__375 clknet_1_1__leaf__02752_ vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__inv_2
XFILLER_124_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10365_ _03246_ vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__clkbuf_1
X_13153_ _05877_ _05884_ _05909_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__a21oi_1
XFILLER_83_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _04850_ _04854_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__and2b_1
XFILLER_112_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17961_ rbzero.pov.spi_buffer\[34\] rbzero.pov.ready_buffer\[34\] _02175_ vssd1 vssd1
+ vccd1 vccd1 _02181_ sky130_fd_sc_hd__mux2_1
X_13084_ _05489_ _05838_ _05840_ _05807_ _05817_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__o2111a_1
XFILLER_69_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10296_ _03072_ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__clkbuf_4
XFILLER_152_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16912_ _09517_ _09518_ _08509_ vssd1 vssd1 vccd1 vccd1 _09519_ sky130_fd_sc_hd__a21oi_1
X_12035_ _04792_ net35 vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__nor2_1
X_19700_ clknet_leaf_73_i_clk _00631_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17892_ rbzero.pov.spi_buffer\[1\] rbzero.pov.ready_buffer\[1\] _02143_ vssd1 vssd1
+ vccd1 vccd1 _02145_ sky130_fd_sc_hd__mux2_1
XFILLER_77_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16843_ _09448_ _09449_ vssd1 vssd1 vccd1 vccd1 _09450_ sky130_fd_sc_hd__xnor2_1
X_19631_ clknet_leaf_53_i_clk _00562_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19562_ clknet_leaf_36_i_clk _00493_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16774_ _09046_ _09381_ vssd1 vssd1 vccd1 vccd1 _09382_ sky130_fd_sc_hd__or2_1
X_13986_ _05318_ _06663_ _06667_ _05373_ _06629_ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__a221oi_2
XFILLER_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18513_ rbzero.pov.spi_buffer\[26\] rbzero.pov.spi_buffer\[27\] _02466_ vssd1 vssd1
+ vccd1 vccd1 _02474_ sky130_fd_sc_hd__mux2_1
X_15725_ _08273_ _08274_ vssd1 vssd1 vccd1 vccd1 _08408_ sky130_fd_sc_hd__and2_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12937_ _05499_ _05688_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19493_ clknet_leaf_46_i_clk _00439_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15656_ _07097_ _07332_ vssd1 vssd1 vccd1 vccd1 _08339_ sky130_fd_sc_hd__or2_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _05623_ _05624_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__or2_1
XFILLER_15_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _07216_ _07294_ vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__xnor2_1
X_18375_ rbzero.pov.spi_counter\[5\] _02426_ _02415_ vssd1 vssd1 vccd1 vccd1 _02429_
+ sky130_fd_sc_hd__a21boi_1
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11819_ gpout2.clk_div\[1\] _04577_ _04570_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__and3_1
X_15587_ _07175_ _04950_ _03493_ _08269_ vssd1 vssd1 vccd1 vccd1 _08271_ sky130_fd_sc_hd__or4_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _05541_ _05542_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__xnor2_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17326_ _01646_ _01647_ _01648_ vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14538_ _07224_ _07225_ vssd1 vssd1 vccd1 vccd1 _07226_ sky130_fd_sc_hd__and2_1
XFILLER_174_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17257_ _04964_ _01527_ _01589_ vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__a21oi_1
X_14469_ _07156_ vssd1 vssd1 vccd1 vccd1 _07157_ sky130_fd_sc_hd__clkbuf_4
X_16208_ _08763_ _08820_ vssd1 vssd1 vccd1 vccd1 _08821_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17188_ rbzero.wall_tracer.trackDistY\[-10\] rbzero.wall_tracer.stepDistY\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__nand2_1
XFILLER_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16139_ _08742_ _08751_ vssd1 vssd1 vccd1 vccd1 _08752_ sky130_fd_sc_hd__nand2_1
XFILLER_115_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19829_ clknet_leaf_20_i_clk _00760_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.vinf
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_110_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19233__8 clknet_1_1__leaf__02754_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__inv_2
XFILLER_20_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_78 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_78/HI o_rgb[5] sky130_fd_sc_hd__conb_1
XFILLER_181_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_89 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_89/HI o_rgb[20] sky130_fd_sc_hd__conb_1
XFILLER_165_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20466_ net146 _01397_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20397_ net457 _01328_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10150_ _03133_ vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10081_ _03097_ vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__clkbuf_1
XFILLER_102_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13840_ _06196_ _06591_ _06596_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__or3_2
XFILLER_62_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13771_ _06526_ _06527_ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__nor2_1
X_10983_ _03636_ _03719_ _03687_ _03535_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__or4_1
XFILLER_28_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15510_ _07269_ _07959_ _08193_ vssd1 vssd1 vccd1 vccd1 _08194_ sky130_fd_sc_hd__or3b_1
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12722_ _05478_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__clkbuf_4
X_16490_ _07984_ _08191_ vssd1 vssd1 vccd1 vccd1 _09100_ sky130_fd_sc_hd__nor2_1
XFILLER_31_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15441_ _08008_ _08117_ _08124_ vssd1 vssd1 vccd1 vccd1 _08126_ sky130_fd_sc_hd__nand3_1
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12653_ _05274_ _05338_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__nor2_2
XFILLER_30_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11604_ rbzero.row_render.wall\[1\] _03997_ _04385_ vssd1 vssd1 vccd1 vccd1 _04386_
+ sky130_fd_sc_hd__and3_1
X_18160_ rbzero.spi_registers.new_mapd\[14\] _02290_ _02297_ _02275_ vssd1 vssd1 vccd1
+ vccd1 _00765_ sky130_fd_sc_hd__o211a_1
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15372_ _07931_ _07934_ _08056_ vssd1 vssd1 vccd1 vccd1 _08058_ sky130_fd_sc_hd__nand3_1
X_12584_ _05201_ _05305_ _05302_ _05306_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__or4_1
XFILLER_196_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17111_ _09709_ _09715_ rbzero.wall_tracer.trackDistX\[9\] _08508_ vssd1 vssd1 vccd1
+ vccd1 _00558_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_50_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14323_ _06866_ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__clkbuf_4
X_11535_ rbzero.tex_b0\[59\] rbzero.tex_b0\[58\] _03732_ vssd1 vssd1 vccd1 vccd1 _04317_
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18091_ _02250_ vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17042_ _09548_ _09551_ _09645_ vssd1 vssd1 vccd1 vccd1 _09647_ sky130_fd_sc_hd__nor3_1
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14254_ rbzero.debug_overlay.playerY\[-5\] vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__inv_2
X_11466_ rbzero.tex_g1\[29\] rbzero.tex_g1\[28\] _04247_ vssd1 vssd1 vccd1 vccd1 _04249_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__02731_ _02731_ vssd1 vssd1 vccd1 vccd1 clknet_0__02731_ sky130_fd_sc_hd__clkbuf_16
X_13205_ _05471_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__inv_2
X_10417_ _03273_ vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__clkbuf_1
X_11397_ rbzero.tex_g0\[9\] rbzero.tex_g0\[8\] _03662_ vssd1 vssd1 vccd1 vccd1 _04181_
+ sky130_fd_sc_hd__mux2_1
X_14185_ _06872_ vssd1 vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__clkbuf_4
XFILLER_125_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13136_ _05533_ _05645_ _05892_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__a21boi_1
X_18934__118 clknet_1_1__leaf__02725_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__inv_2
X_10348_ _03237_ vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10279_ _03201_ vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17944_ rbzero.pov.spi_buffer\[26\] rbzero.pov.ready_buffer\[26\] _02164_ vssd1 vssd1
+ vccd1 vccd1 _02172_ sky130_fd_sc_hd__mux2_1
X_13067_ _05819_ _05823_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__or2_1
X_12018_ net34 _04790_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__nor2_1
XFILLER_39_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17875_ rbzero.spi_registers.spi_counter\[3\] _02102_ _02103_ _02132_ vssd1 vssd1
+ vccd1 vccd1 _00645_ sky130_fd_sc_hd__o211a_1
XFILLER_66_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19614_ clknet_leaf_60_i_clk _00545_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16826_ _08862_ _08071_ vssd1 vssd1 vccd1 vccd1 _09433_ sky130_fd_sc_hd__nor2_1
XFILLER_65_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16757_ _09021_ _09039_ vssd1 vssd1 vccd1 vccd1 _09365_ sky130_fd_sc_hd__nor2_1
XFILLER_4_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19545_ clknet_leaf_37_i_clk _00476_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13969_ _05270_ _06636_ _06637_ _06716_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__a31o_4
XFILLER_0_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15708_ _04841_ rbzero.wall_tracer.stepDistX\[8\] _08141_ _08390_ vssd1 vssd1 vccd1
+ vccd1 _08391_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16688_ _09295_ _09296_ vssd1 vssd1 vccd1 vccd1 _09297_ sky130_fd_sc_hd__nor2_1
X_19476_ clknet_leaf_54_i_clk _00422_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15639_ _08221_ _08288_ vssd1 vssd1 vccd1 vccd1 _08322_ sky130_fd_sc_hd__nand2_1
XFILLER_62_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18358_ rbzero.pov.spi_counter\[0\] _02414_ _02416_ vssd1 vssd1 vccd1 vccd1 _00844_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_147_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17309_ rbzero.wall_tracer.trackDistY\[7\] rbzero.wall_tracer.stepDistY\[7\] vssd1
+ vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__nor2_1
XFILLER_175_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18289_ _02370_ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__inv_2
XFILLER_175_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20320_ net380 _01251_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20251_ net311 _01182_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20182_ net242 _01113_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[29\] sky130_fd_sc_hd__dfxtp_1
X_09993_ rbzero.tex_r0\[4\] rbzero.tex_r0\[3\] _03050_ vssd1 vssd1 vccd1 vccd1 _03051_
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11320_ rbzero.debug_overlay.vplaneX\[0\] _04079_ _04099_ _04104_ vssd1 vssd1 vccd1
+ vccd1 _04105_ sky130_fd_sc_hd__a211o_1
X_20518_ clknet_leaf_27_i_clk _01449_ vssd1 vssd1 vccd1 vccd1 gpout1.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11251_ gpout0.hpos\[7\] _03512_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__nor2_1
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20449_ net129 _01380_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10202_ rbzero.tex_g0\[33\] rbzero.tex_g0\[32\] _03155_ vssd1 vssd1 vccd1 vccd1 _03161_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11182_ _03960_ _03962_ _03964_ _03966_ _03721_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__o221a_1
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10133_ _03124_ vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15990_ _08335_ _08350_ _08348_ vssd1 vssd1 vccd1 vccd1 _08604_ sky130_fd_sc_hd__a21o_1
X_14941_ _07621_ _07627_ _07628_ vssd1 vssd1 vccd1 vccd1 _07629_ sky130_fd_sc_hd__a21oi_1
X_10064_ _03088_ vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_130_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17660_ _01933_ _01934_ _01935_ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__and3_1
XFILLER_75_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14872_ _07552_ _07558_ _07559_ vssd1 vssd1 vccd1 vccd1 _07560_ sky130_fd_sc_hd__a21oi_1
X_19029__204 clknet_1_0__leaf__02734_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__inv_2
XFILLER_78_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16611_ _09214_ _09219_ vssd1 vssd1 vccd1 vccd1 _09220_ sky130_fd_sc_hd__xnor2_1
XFILLER_85_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13823_ _06198_ _06201_ _06578_ _06579_ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__a31o_1
XFILLER_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17591_ _01862_ _01870_ _01874_ _01876_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__a31o_1
XFILLER_29_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16542_ _09150_ _09151_ vssd1 vssd1 vccd1 vccd1 _09152_ sky130_fd_sc_hd__nand2_1
X_19330_ _02759_ _02814_ _02815_ _02319_ rbzero.texV\[0\] vssd1 vssd1 vccd1 vccd1
+ _01417_ sky130_fd_sc_hd__a32o_1
X_13754_ _06500_ _06506_ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__xnor2_1
X_10966_ _03659_ _03751_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__or2_1
XFILLER_188_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19261_ _02758_ vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12705_ _05461_ _05434_ _05376_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__mux2_1
X_16473_ _08960_ _08965_ vssd1 vssd1 vccd1 vccd1 _09084_ sky130_fd_sc_hd__nand2_1
X_13685_ _06103_ _06156_ vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__nor2_1
XFILLER_188_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10897_ _03596_ _03682_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__xnor2_2
X_18212_ _02323_ _02328_ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__and2_1
X_15424_ _08107_ _08108_ _07980_ _07979_ _07860_ vssd1 vssd1 vccd1 vccd1 _08109_ sky130_fd_sc_hd__o32a_1
XFILLER_148_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12636_ _05338_ _05383_ _05386_ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__and3_1
XFILLER_157_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18143_ rbzero.spi_registers.new_vinf _02278_ _02283_ _02284_ _02285_ vssd1 vssd1
+ vccd1 vccd1 _00760_ sky130_fd_sc_hd__o311a_1
XFILLER_200_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15355_ _07850_ _07917_ _07916_ vssd1 vssd1 vccd1 vccd1 _08041_ sky130_fd_sc_hd__a21oi_1
X_12567_ _05313_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__clkbuf_4
XFILLER_129_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14306_ _06979_ _06993_ vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__nor2_1
X_11518_ rbzero.tex_g1\[46\] _03733_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__and2_1
X_18074_ rbzero.spi_registers.spi_buffer\[13\] rbzero.spi_registers.spi_buffer\[12\]
+ _02226_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__mux2_1
X_15286_ _06979_ vssd1 vssd1 vccd1 vccd1 _07972_ sky130_fd_sc_hd__buf_2
XFILLER_184_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12498_ _05223_ _05254_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__nor2_1
X_19075__246 clknet_1_1__leaf__02738_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__inv_2
X_17025_ _09601_ _09602_ vssd1 vssd1 vccd1 vccd1 _09630_ sky130_fd_sc_hd__or2_1
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14237_ rbzero.debug_overlay.playerY\[-6\] _06924_ _04928_ vssd1 vssd1 vccd1 vccd1
+ _06925_ sky130_fd_sc_hd__mux2_1
X_11449_ _03896_ _04230_ _04232_ _03522_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__a211o_1
XFILLER_125_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14168_ rbzero.wall_tracer.visualWallDist\[1\] _06855_ vssd1 vssd1 vccd1 vccd1 _06856_
+ sky130_fd_sc_hd__nand2_1
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _05625_ _05617_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__and2b_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18976_ clknet_1_1__leaf__02440_ vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__buf_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14099_ rbzero.wall_tracer.trackDistX\[9\] _05004_ _06812_ _06813_ _06783_ vssd1
+ vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__a221o_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17927_ rbzero.pov.spi_buffer\[18\] rbzero.pov.ready_buffer\[18\] _02153_ vssd1 vssd1
+ vccd1 vccd1 _02163_ sky130_fd_sc_hd__mux2_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17858_ rbzero.spi_registers.spi_counter\[4\] _01659_ _02118_ vssd1 vssd1 vccd1 vccd1
+ _02119_ sky130_fd_sc_hd__o21ai_1
XFILLER_82_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18443__82 clknet_1_1__leaf__02439_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__inv_2
X_16809_ rbzero.wall_tracer.trackDistX\[6\] rbzero.wall_tracer.stepDistX\[6\] vssd1
+ vssd1 vccd1 vccd1 _09417_ sky130_fd_sc_hd__nor2_1
X_17789_ _02000_ rbzero.debug_overlay.vplaneX\[-2\] vssd1 vssd1 vccd1 vccd1 _02055_
+ sky130_fd_sc_hd__nand2_1
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19528_ clknet_leaf_66_i_clk _00000_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19459_ clknet_leaf_64_i_clk _00405_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_201_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20303_ net363 _01234_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20234_ net294 _01165_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20165_ net225 _01096_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[12\] sky130_fd_sc_hd__dfxtp_1
X_09976_ rbzero.tex_r0\[12\] rbzero.tex_r0\[11\] _03039_ vssd1 vssd1 vccd1 vccd1 _03042_
+ sky130_fd_sc_hd__mux2_1
XFILLER_118_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20096_ clknet_leaf_90_i_clk _01027_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10820_ _03605_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__buf_4
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10751_ net41 vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__buf_4
XFILLER_52_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13470_ _06224_ _06226_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__nor2_1
XFILLER_125_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10682_ _03471_ _03472_ _03475_ _03476_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__or4_1
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12421_ _05163_ _05177_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__xor2_2
XFILLER_185_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15140_ _07824_ _07827_ vssd1 vssd1 vccd1 vccd1 _07828_ sky130_fd_sc_hd__nor2_1
XFILLER_154_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12352_ rbzero.wall_tracer.visualWallDist\[-8\] rbzero.wall_tracer.rcp_sel\[2\] _05072_
+ _05108_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__o211a_1
XFILLER_181_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11303_ rbzero.debug_overlay.facingY\[0\] _04079_ _04081_ rbzero.debug_overlay.facingY\[-9\]
+ _04087_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__a221o_1
X_15071_ _07755_ _07758_ vssd1 vssd1 vccd1 vccd1 _07759_ sky130_fd_sc_hd__nand2_1
X_12283_ rbzero.debug_overlay.facingX\[-9\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__nand2_2
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14022_ _06675_ _05390_ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__nor2_1
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11234_ _03461_ _02901_ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__nor2_1
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18830_ rbzero.pov.ready_buffer\[18\] _02666_ _02677_ _02675_ vssd1 vssd1 vccd1 vccd1
+ _01055_ sky130_fd_sc_hd__a211o_1
XFILLER_106_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11165_ rbzero.tex_r1\[37\] _03659_ _03767_ _03606_ vssd1 vssd1 vccd1 vccd1 _03950_
+ sky130_fd_sc_hd__a31o_1
XFILLER_136_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10116_ _03115_ vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18761_ _02637_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__clkbuf_2
XFILLER_49_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11096_ gpout0.vpos\[4\] rbzero.map_overlay.i_othery\[1\] vssd1 vssd1 vccd1 vccd1
+ _03882_ sky130_fd_sc_hd__xor2_1
X_15973_ _08578_ _08580_ _08579_ vssd1 vssd1 vccd1 vccd1 _08588_ sky130_fd_sc_hd__a21boi_1
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14924_ _07576_ _07608_ vssd1 vssd1 vccd1 vccd1 _07612_ sky130_fd_sc_hd__nand2_1
X_10047_ _03079_ vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__clkbuf_1
X_17712_ rbzero.wall_tracer.rayAddendX\[0\] _01983_ _03509_ vssd1 vssd1 vccd1 vccd1
+ _01984_ sky130_fd_sc_hd__mux2_1
XFILLER_48_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18692_ _02583_ rbzero.pov.ready_buffer\[44\] _02535_ vssd1 vssd1 vccd1 vccd1 _02584_
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14855_ _06873_ _07530_ _07539_ _07541_ _07542_ vssd1 vssd1 vccd1 vccd1 _07543_ sky130_fd_sc_hd__o41a_1
X_17643_ rbzero.debug_overlay.vplaneX\[-7\] rbzero.wall_tracer.rayAddendX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__nor2_1
XFILLER_1_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13806_ _06432_ _06335_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__and2_1
X_17574_ _01859_ _01860_ _01845_ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__o21ai_1
X_14786_ _07425_ _07426_ _07473_ vssd1 vssd1 vccd1 vccd1 _07474_ sky130_fd_sc_hd__o21a_1
X_11998_ _04750_ net62 _04771_ net31 vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__o211a_1
XFILLER_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16525_ _09009_ _09133_ _09008_ vssd1 vssd1 vccd1 vccd1 _09135_ sky130_fd_sc_hd__o21bai_1
X_19313_ rbzero.traced_texa\[-2\] rbzero.texV\[-2\] vssd1 vssd1 vccd1 vccd1 _02801_
+ sky130_fd_sc_hd__nand2_1
XFILLER_95_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13737_ _06492_ _06493_ vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__nor2_1
XFILLER_95_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10949_ _03726_ _03728_ _03731_ _03734_ _03674_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__o221a_1
XFILLER_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16456_ _08882_ _08942_ _08940_ vssd1 vssd1 vccd1 vccd1 _09067_ sky130_fd_sc_hd__a21oi_1
X_13668_ _06397_ _06423_ _06424_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__a21o_1
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15407_ _08068_ _08091_ vssd1 vssd1 vccd1 vccd1 _08092_ sky130_fd_sc_hd__xnor2_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12619_ _05375_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__clkbuf_4
X_16387_ _08996_ _08997_ vssd1 vssd1 vccd1 vccd1 _08998_ sky130_fd_sc_hd__nor2_1
XFILLER_31_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13599_ _06342_ _06351_ _06353_ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__and3_1
XFILLER_145_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18126_ rbzero.map_overlay.i_othery\[1\] _02268_ vssd1 vssd1 vccd1 vccd1 _02273_
+ sky130_fd_sc_hd__or2_1
X_15338_ _07673_ _07173_ _07901_ _07899_ vssd1 vssd1 vccd1 vccd1 _08024_ sky130_fd_sc_hd__a31oi_1
XFILLER_129_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18057_ _02232_ vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15269_ _07843_ _07954_ vssd1 vssd1 vccd1 vccd1 _07955_ sky130_fd_sc_hd__nor2_1
X_17008_ _09611_ _09612_ vssd1 vssd1 vccd1 vccd1 _09614_ sky130_fd_sc_hd__and2_1
XFILLER_126_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09830_ _02963_ vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09761_ _02927_ vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18986__166 clknet_1_0__leaf__02729_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__inv_2
XFILLER_199_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19058__230 clknet_1_1__leaf__02737_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__inv_2
XFILLER_109_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20217_ net277 _01148_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20148_ clknet_leaf_13_i_clk _01079_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[6\] sky130_fd_sc_hd__dfxtp_4
X_09959_ rbzero.tex_r0\[20\] rbzero.tex_r0\[19\] _03028_ vssd1 vssd1 vccd1 vccd1 _03033_
+ sky130_fd_sc_hd__mux2_1
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12970_ _05691_ _05692_ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__xnor2_1
X_20079_ clknet_leaf_7_i_clk _01010_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_46_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ _04507_ _04508_ _03520_ _03515_ net21 _04670_ vssd1 vssd1 vccd1 vccd1 _04696_
+ sky130_fd_sc_hd__mux4_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _07318_ _07326_ _07327_ vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__a21oi_2
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18422__63 clknet_1_0__leaf__02437_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__inv_2
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ net40 _04626_ _04627_ _03537_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__a22o_1
XFILLER_33_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _03585_ _03586_ _03588_ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__nand3_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _07255_ _07258_ vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__xnor2_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _04552_ net65 _04558_ _04559_ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__a211o_1
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16310_ _08920_ _08921_ vssd1 vssd1 vccd1 vccd1 _08922_ sky130_fd_sc_hd__and2_1
XFILLER_158_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13522_ _06140_ _06191_ vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__and2_1
XFILLER_198_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10734_ gpout0.vpos\[6\] vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__clkbuf_4
X_17290_ _01616_ _01617_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__nand2_1
XFILLER_201_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16241_ _08851_ _08852_ vssd1 vssd1 vccd1 vccd1 _08853_ sky130_fd_sc_hd__nor2_1
X_13453_ _06208_ _06209_ vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__nor2_1
XFILLER_201_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10665_ gpout0.hpos\[5\] vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__buf_4
XFILLER_185_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12404_ _03488_ _05078_ _05160_ _05080_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__o31a_2
X_16172_ _08783_ _08784_ vssd1 vssd1 vccd1 vccd1 _08785_ sky130_fd_sc_hd__nand2_1
XFILLER_167_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13384_ _06073_ _06075_ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__and2_1
XFILLER_139_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10596_ _03390_ _03358_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__or2_1
XFILLER_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15123_ _07808_ _07809_ vssd1 vssd1 vccd1 vccd1 _07811_ sky130_fd_sc_hd__or2_1
X_12335_ _03479_ _04905_ _04906_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__and3_1
XFILLER_86_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19931_ net160 _00862_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[11\] sky130_fd_sc_hd__dfxtp_1
X_15054_ _07646_ _07198_ vssd1 vssd1 vccd1 vccd1 _07742_ sky130_fd_sc_hd__nor2_1
XFILLER_126_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12266_ rbzero.wall_tracer.mapY\[9\] _04923_ _05023_ vssd1 vssd1 vccd1 vccd1 _05024_
+ sky130_fd_sc_hd__a21o_1
X_14005_ _06708_ _06723_ _06664_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__mux2_1
X_11217_ _03996_ _03999_ _04000_ _04001_ _03764_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__a221o_1
XFILLER_141_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19862_ clknet_leaf_23_i_clk _00793_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 o_tex_out0 sky130_fd_sc_hd__buf_2
X_12197_ rbzero.wall_tracer.trackDistY\[5\] vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__inv_2
XFILLER_68_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_1_1_0_i_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_150_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18813_ _01967_ _02666_ vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__nor2_1
XFILLER_68_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11148_ rbzero.tex_r1\[60\] _03920_ _03925_ _03932_ vssd1 vssd1 vccd1 vccd1 _03933_
+ sky130_fd_sc_hd__a31o_1
XFILLER_1_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19793_ clknet_leaf_18_i_clk _00724_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18744_ _02623_ vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__clkbuf_1
X_11079_ _02900_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__clkinv_4
X_15956_ _08570_ _08571_ _08572_ vssd1 vssd1 vccd1 vccd1 _08573_ sky130_fd_sc_hd__nor3_1
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14907_ _07533_ _07577_ _07578_ vssd1 vssd1 vccd1 vccd1 _07595_ sky130_fd_sc_hd__a21o_1
XFILLER_37_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18675_ rbzero.debug_overlay.playerX\[3\] _02566_ vssd1 vssd1 vccd1 vccd1 _02570_
+ sky130_fd_sc_hd__or2_1
X_15887_ _08509_ vssd1 vssd1 vccd1 vccd1 _08512_ sky130_fd_sc_hd__buf_4
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17626_ rbzero.debug_overlay.playerY\[3\] _01905_ _09620_ vssd1 vssd1 vccd1 vccd1
+ _01906_ sky130_fd_sc_hd__mux2_1
X_14838_ _07479_ _07525_ vssd1 vssd1 vccd1 vccd1 _07526_ sky130_fd_sc_hd__and2_1
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17557_ _01784_ _04109_ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__or2_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14769_ _07448_ _07454_ vssd1 vssd1 vccd1 vccd1 _07457_ sky130_fd_sc_hd__xor2_1
X_16508_ _09112_ _09117_ vssd1 vssd1 vccd1 vccd1 _09118_ sky130_fd_sc_hd__and2_1
X_17488_ _01764_ _01766_ _01765_ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__a21bo_1
XFILLER_32_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16439_ _07877_ _09049_ vssd1 vssd1 vccd1 vccd1 _09050_ sky130_fd_sc_hd__or2_1
XFILLER_192_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18109_ _02261_ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__buf_4
XFILLER_117_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20002_ clknet_leaf_93_i_clk _00933_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_09813_ rbzero.tex_r1\[23\] rbzero.tex_r1\[24\] _02954_ vssd1 vssd1 vccd1 vccd1 _02955_
+ sky130_fd_sc_hd__mux2_1
XFILLER_119_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09744_ _02918_ vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_i_clk clknet_2_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10450_ _03290_ vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10381_ rbzero.tex_b1\[11\] rbzero.tex_b1\[12\] _03254_ vssd1 vssd1 vccd1 vccd1 _03255_
+ sky130_fd_sc_hd__mux2_1
XFILLER_109_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12120_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[10\] vssd1
+ vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__or2_1
XFILLER_108_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12051_ _04801_ _04820_ _04823_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__o21ba_2
XFILLER_123_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11002_ rbzero.row_render.size\[4\] _03463_ _03782_ rbzero.row_render.size\[5\] _03787_
+ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__a221o_1
XFILLER_172_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15810_ rbzero.traced_texa\[-7\] _08457_ _08459_ rbzero.wall_tracer.visualWallDist\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__a22o_1
X_16790_ _09245_ _09292_ _09397_ vssd1 vssd1 vccd1 vccd1 _09398_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15741_ _08320_ _08423_ vssd1 vssd1 vccd1 vccd1 _08424_ sky130_fd_sc_hd__xnor2_1
XFILLER_133_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ _05473_ _05551_ _05610_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__mux2_1
X_18969__150 clknet_1_1__leaf__02728_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__inv_2
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11904_ net24 _04670_ net25 vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__a21oi_1
X_15672_ _08323_ _08354_ vssd1 vssd1 vccd1 vccd1 _08355_ sky130_fd_sc_hd__xnor2_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18460_ _02446_ vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__clkbuf_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _05631_ _05640_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__nor2_1
XFILLER_46_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _07234_ _07236_ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__xnor2_1
X_17411_ _01704_ _01708_ _01709_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__o21ai_1
XFILLER_73_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _04562_ _04610_ _04611_ net66 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__o22a_2
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _01662_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__clkbuf_4
X_14554_ _07237_ _07241_ vssd1 vssd1 vccd1 vccd1 _07242_ sky130_fd_sc_hd__xnor2_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _04542_ _04543_ net6 vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__mux2_1
XFILLER_186_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _06122_ _06035_ _06128_ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__or3_1
X_10717_ _03464_ _03461_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__nor2_1
X_17273_ rbzero.wall_tracer.trackDistY\[2\] rbzero.wall_tracer.stepDistY\[2\] vssd1
+ vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__or2_1
X_14485_ _07171_ _07172_ _04841_ rbzero.wall_tracer.stepDistX\[4\] vssd1 vssd1 vccd1
+ vccd1 _07173_ sky130_fd_sc_hd__o2bb2a_4
X_11697_ _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__inv_2
XFILLER_201_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16224_ rbzero.wall_tracer.trackDistX\[1\] rbzero.wall_tracer.stepDistX\[1\] vssd1
+ vssd1 vccd1 vccd1 _08837_ sky130_fd_sc_hd__or2_1
X_13436_ _05997_ _06095_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__nand2_1
X_10648_ _03436_ _03439_ _03440_ _03443_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__or4_1
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16155_ _07012_ _07878_ vssd1 vssd1 vccd1 vccd1 _08768_ sky130_fd_sc_hd__nor2_1
XFILLER_154_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13367_ _06121_ _06123_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__or2_1
X_10579_ rbzero.map_rom.a6 vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__clkinv_2
XFILLER_177_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15106_ _07782_ _07792_ vssd1 vssd1 vccd1 vccd1 _07794_ sky130_fd_sc_hd__or2_1
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12318_ _05073_ _05074_ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__xnor2_2
XFILLER_182_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16086_ _08697_ _08698_ vssd1 vssd1 vccd1 vccd1 _08700_ sky130_fd_sc_hd__nand2_1
X_13298_ _06002_ _06034_ _06054_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__a21oi_4
XFILLER_170_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15037_ _07125_ _07705_ _07723_ vssd1 vssd1 vccd1 vccd1 _07725_ sky130_fd_sc_hd__nand3_1
X_19914_ clknet_leaf_0_i_clk _00845_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12249_ rbzero.wall_tracer.mapY\[7\] _04923_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19845_ clknet_leaf_18_i_clk _00776_ vssd1 vssd1 vccd1 vccd1 rbzero.mapdyw\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_95_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19776_ clknet_leaf_5_i_clk _00707_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_16988_ _09592_ _09593_ vssd1 vssd1 vccd1 vccd1 _09594_ sky130_fd_sc_hd__nand2_1
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18727_ rbzero.debug_overlay.playerY\[0\] _02588_ _02609_ _02586_ vssd1 vssd1 vccd1
+ vccd1 _01020_ sky130_fd_sc_hd__o211a_1
XFILLER_114_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15939_ _08555_ _08556_ _08557_ vssd1 vssd1 vccd1 vccd1 _08558_ sky130_fd_sc_hd__or3_1
XFILLER_97_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18658_ _07034_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__inv_2
XFILLER_24_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17609_ rbzero.wall_tracer.rayAddendY\[10\] _01892_ _03509_ vssd1 vssd1 vccd1 vccd1
+ _01893_ sky130_fd_sc_hd__mux2_1
XFILLER_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18401__44 clknet_1_1__leaf__02435_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__inv_2
X_18589_ rbzero.pov.spi_buffer\[62\] rbzero.pov.spi_buffer\[63\] _02510_ vssd1 vssd1
+ vccd1 vccd1 _02514_ sky130_fd_sc_hd__mux2_1
XFILLER_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20482_ clknet_leaf_61_i_clk _01413_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09727_ _02908_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__buf_4
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _03611_ _04400_ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__or2_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11551_ rbzero.tex_b0\[35\] _04155_ _04156_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__and3_1
XFILLER_184_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10502_ rbzero.tex_b0\[18\] rbzero.tex_b0\[17\] _03313_ vssd1 vssd1 vccd1 vccd1 _03318_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14270_ _06956_ _06957_ vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__and2_1
XFILLER_109_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11482_ rbzero.tex_g1\[7\] rbzero.tex_g1\[6\] _04247_ vssd1 vssd1 vccd1 vccd1 _04265_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13221_ _05936_ _05939_ _05977_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__a21oi_4
XFILLER_171_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10433_ rbzero.tex_b0\[51\] rbzero.tex_b0\[50\] _03280_ vssd1 vssd1 vccd1 vccd1 _03282_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13152_ _05636_ _05885_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__nor2_1
XFILLER_109_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10364_ rbzero.tex_b1\[19\] rbzero.tex_b1\[20\] _03243_ vssd1 vssd1 vccd1 vccd1 _03246_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ _04849_ _04856_ _04857_ _04864_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__or4bb_1
XFILLER_124_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17960_ _02180_ vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__clkbuf_1
X_13083_ _05516_ _05551_ _05549_ _05697_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10295_ _03209_ vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__clkbuf_1
X_16911_ _09408_ _09415_ vssd1 vssd1 vccd1 vccd1 _09518_ sky130_fd_sc_hd__nand2_1
X_12034_ _04507_ _04508_ _03520_ _03515_ _04790_ net35 vssd1 vssd1 vccd1 vccd1 _04807_
+ sky130_fd_sc_hd__mux4_1
XFILLER_77_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17891_ _02144_ vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19630_ clknet_leaf_53_i_clk _00561_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
X_16842_ _08899_ _09110_ vssd1 vssd1 vccd1 vccd1 _09449_ sky130_fd_sc_hd__nor2_1
XFILLER_19_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19561_ clknet_leaf_63_i_clk _00492_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16773_ _07992_ _09379_ vssd1 vssd1 vccd1 vccd1 _09381_ sky130_fd_sc_hd__or2b_1
XFILLER_19_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13985_ _06701_ _06730_ _05310_ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__mux2_1
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18512_ _02473_ vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__clkbuf_1
X_15724_ _08395_ _08406_ vssd1 vssd1 vccd1 vccd1 _08407_ sky130_fd_sc_hd__xnor2_2
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12936_ _05654_ _05690_ _05691_ _05692_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__o2bb2a_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19492_ clknet_leaf_39_i_clk _00438_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15655_ _07984_ _07270_ _08226_ vssd1 vssd1 vccd1 vccd1 _08338_ sky130_fd_sc_hd__or3_1
X_12867_ _05619_ _05580_ _05622_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__and3_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14606_ _07141_ _07148_ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__nor2_1
X_11818_ _04532_ _04571_ _04565_ _04570_ _04594_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__a41o_1
X_18374_ _02428_ vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15586_ _04950_ _08269_ _06860_ rbzero.wall_tracer.visualWallDist\[-10\] vssd1 vssd1
+ vccd1 vccd1 _08270_ sky130_fd_sc_hd__and4bb_2
X_12798_ _05544_ _05554_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__xor2_2
XFILLER_15_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17325_ _01640_ _01642_ _01641_ vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__a21bo_1
X_14537_ _07078_ _06933_ _07221_ _07223_ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__a2bb2o_1
X_11749_ net7 vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__inv_2
XFILLER_187_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14468_ _06787_ _06855_ vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__nand2_2
X_17256_ _08485_ _01587_ _01588_ _08584_ _01522_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__o311a_1
X_16207_ _08817_ _08819_ vssd1 vssd1 vccd1 vccd1 _08820_ sky130_fd_sc_hd__xor2_1
X_13419_ _06166_ _06175_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__or2_1
X_17187_ rbzero.wall_tracer.trackDistY\[-10\] rbzero.wall_tracer.stepDistY\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__or2_1
XFILLER_143_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14399_ _06859_ rbzero.wall_tracer.stepDistY\[-2\] _04838_ vssd1 vssd1 vccd1 vccd1
+ _07087_ sky130_fd_sc_hd__o21ai_1
X_16138_ _08749_ _08750_ vssd1 vssd1 vccd1 vccd1 _08751_ sky130_fd_sc_hd__and2_1
XFILLER_6_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16069_ _07185_ _07199_ vssd1 vssd1 vccd1 vccd1 _08683_ sky130_fd_sc_hd__nand2_1
XFILLER_88_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19828_ clknet_leaf_13_i_clk _00759_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19759_ clknet_leaf_87_i_clk _00690_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtop_ew_algofoogle_79 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_79/HI o_rgb[8] sky130_fd_sc_hd__conb_1
X_20465_ net145 _01396_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20396_ net456 _01327_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10080_ rbzero.tex_g1\[26\] rbzero.tex_g1\[27\] _03095_ vssd1 vssd1 vccd1 vccd1 _03097_
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13770_ _06525_ _06514_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__and2b_1
X_10982_ _03767_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_40_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12721_ _05454_ _05455_ _05457_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__or3b_1
XFILLER_74_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15440_ _08008_ _08117_ _08124_ vssd1 vssd1 vccd1 vccd1 _08125_ sky130_fd_sc_hd__a21o_1
Xclkbuf_2_0_0_i_clk clknet_1_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_70_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19224__380 clknet_1_1__leaf__02753_ vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__inv_2
X_12652_ _05212_ _05238_ _05311_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__mux2_1
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11603_ _04179_ _04192_ _03768_ _03631_ rbzero.row_render.side vssd1 vssd1 vccd1
+ vccd1 _04385_ sky130_fd_sc_hd__a311o_1
XFILLER_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15371_ _07931_ _07934_ _08056_ vssd1 vssd1 vccd1 vccd1 _08057_ sky130_fd_sc_hd__a21o_1
X_12583_ _05244_ _05276_ _05297_ _05231_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__a31o_1
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_55_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_17110_ _09713_ _09714_ _08507_ vssd1 vssd1 vccd1 vccd1 _09715_ sky130_fd_sc_hd__o21a_1
X_14322_ _06941_ _06995_ _07009_ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__a21bo_1
XFILLER_12_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11534_ rbzero.tex_b0\[57\] rbzero.tex_b0\[56\] _04189_ vssd1 vssd1 vccd1 vccd1 _04316_
+ sky130_fd_sc_hd__mux2_1
XFILLER_129_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18090_ net43 rbzero.spi_registers.mosi_buffer\[0\] _03337_ vssd1 vssd1 vccd1 vccd1
+ _02250_ sky130_fd_sc_hd__mux2_1
XFILLER_184_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17041_ _09548_ _09551_ _09645_ vssd1 vssd1 vccd1 vccd1 _09646_ sky130_fd_sc_hd__o21a_1
XFILLER_128_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14253_ _06921_ _06933_ _06940_ _06920_ vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__o31ai_4
X_11465_ rbzero.tex_g1\[31\] rbzero.tex_g1\[30\] _04247_ vssd1 vssd1 vccd1 vccd1 _04248_
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__02730_ _02730_ vssd1 vssd1 vccd1 vccd1 clknet_0__02730_ sky130_fd_sc_hd__clkbuf_16
XFILLER_171_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13204_ _05912_ _05917_ _05960_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__o21ai_1
X_10416_ rbzero.tex_b0\[59\] rbzero.tex_b0\[58\] _03269_ vssd1 vssd1 vccd1 vccd1 _03273_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14184_ _06871_ vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__clkbuf_4
X_11396_ _03612_ _04176_ _04178_ _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__o211a_1
XFILLER_152_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13135_ _05603_ _05644_ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__or2b_1
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10347_ rbzero.tex_b1\[27\] rbzero.tex_b1\[28\] _03232_ vssd1 vssd1 vccd1 vccd1 _03237_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ _02171_ vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__clkbuf_1
X_13066_ _05819_ _05821_ _05822_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__nor3_1
X_10278_ rbzero.tex_b1\[60\] rbzero.tex_b1\[61\] _03199_ vssd1 vssd1 vccd1 vccd1 _03201_
+ sky130_fd_sc_hd__mux2_1
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12017_ net33 vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__clkbuf_4
XFILLER_94_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17874_ _02122_ _02130_ _02131_ _02123_ vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__a31o_1
XFILLER_38_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19613_ clknet_leaf_60_i_clk _00544_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16825_ _09372_ _09431_ vssd1 vssd1 vccd1 vccd1 _09432_ sky130_fd_sc_hd__nand2_1
XFILLER_65_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19544_ clknet_leaf_41_i_clk _00475_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16756_ _09362_ _09363_ vssd1 vssd1 vccd1 vccd1 _09364_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13968_ _05476_ _06715_ _05272_ vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__a21o_1
XFILLER_59_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15707_ _03493_ rbzero.wall_tracer.stepDistY\[8\] _04950_ vssd1 vssd1 vccd1 vccd1
+ _08390_ sky130_fd_sc_hd__a21oi_1
XFILLER_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12919_ _05658_ _05659_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__xnor2_1
X_19475_ clknet_leaf_49_i_clk _00421_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16687_ _09293_ _09294_ vssd1 vssd1 vccd1 vccd1 _09296_ sky130_fd_sc_hd__and2_1
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13899_ _06603_ _06589_ _06653_ _05271_ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__a211o_1
XFILLER_185_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18426_ clknet_1_0__leaf__02433_ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__buf_1
X_15638_ _08286_ _08287_ vssd1 vssd1 vccd1 vccd1 _08321_ sky130_fd_sc_hd__or2_1
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18357_ rbzero.pov.spi_counter\[0\] _02414_ _02415_ vssd1 vssd1 vccd1 vccd1 _02416_
+ sky130_fd_sc_hd__o21ai_1
X_15569_ _06997_ _08252_ vssd1 vssd1 vccd1 vccd1 _08253_ sky130_fd_sc_hd__nor2_1
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17308_ rbzero.wall_tracer.trackDistY\[6\] _01558_ _01633_ _09416_ vssd1 vssd1 vccd1
+ vccd1 _00577_ sky130_fd_sc_hd__o22a_1
XFILLER_174_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18288_ _02376_ vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__clkbuf_1
XFILLER_163_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17239_ _01566_ _01568_ _01567_ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__a21boi_1
XFILLER_174_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20250_ net310 _01181_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20181_ net241 _01112_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09992_ _02983_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__clkbuf_4
X_19052__225 clknet_1_0__leaf__02736_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__inv_2
XFILLER_170_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19245__19 clknet_1_0__leaf__02755_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__inv_2
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20517_ clknet_leaf_77_i_clk _01448_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_193_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11250_ _03466_ _04034_ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__xnor2_4
XFILLER_107_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20448_ net508 _01379_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10201_ _03160_ vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__clkbuf_1
X_11181_ rbzero.tex_r1\[0\] _03661_ _03936_ _03965_ vssd1 vssd1 vccd1 vccd1 _03966_
+ sky130_fd_sc_hd__a31o_1
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20379_ net439 _01310_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_161_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10132_ rbzero.tex_g1\[1\] rbzero.tex_g1\[2\] _03117_ vssd1 vssd1 vccd1 vccd1 _03124_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18429__69 clknet_1_1__leaf__02438_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__inv_2
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14940_ _07622_ _07626_ vssd1 vssd1 vccd1 vccd1 _07628_ sky130_fd_sc_hd__nor2_1
X_10063_ rbzero.tex_g1\[34\] rbzero.tex_g1\[35\] _03084_ vssd1 vssd1 vccd1 vccd1 _03088_
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14871_ _07553_ _07557_ vssd1 vssd1 vccd1 vccd1 _07559_ sky130_fd_sc_hd__and2b_1
XFILLER_91_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16610_ _09217_ _09218_ vssd1 vssd1 vccd1 vccd1 _09219_ sky130_fd_sc_hd__nor2_1
XFILLER_169_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13822_ _06218_ _06578_ vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__nor2_1
X_17590_ _03339_ _01875_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__nand2_1
XFILLER_91_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16541_ _09042_ _09132_ _09149_ vssd1 vssd1 vccd1 vccd1 _09151_ sky130_fd_sc_hd__nand3_1
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13753_ _06436_ _06469_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__nand2_1
X_10965_ rbzero.tex_r0\[63\] rbzero.tex_r0\[62\] _03662_ vssd1 vssd1 vccd1 vccd1 _03751_
+ sky130_fd_sc_hd__mux2_1
XFILLER_189_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12704_ _05212_ _05215_ _05382_ _05217_ _05349_ _05367_ vssd1 vssd1 vccd1 vccd1 _05461_
+ sky130_fd_sc_hd__mux4_1
X_19260_ _02334_ _02756_ _02757_ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__and3_1
X_13684_ _05527_ _06061_ _06071_ _05862_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__o22ai_1
X_16472_ rbzero.wall_tracer.trackDistX\[3\] rbzero.wall_tracer.stepDistX\[3\] vssd1
+ vssd1 vccd1 vccd1 _09083_ sky130_fd_sc_hd__or2_1
X_10896_ _03681_ _03597_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__nor2_1
X_18211_ rbzero.color_sky\[3\] rbzero.spi_registers.new_sky\[3\] _02320_ vssd1 vssd1
+ vccd1 vccd1 _02328_ sky130_fd_sc_hd__mux2_1
X_15423_ _07281_ vssd1 vssd1 vccd1 vccd1 _08108_ sky130_fd_sc_hd__buf_2
XFILLER_19_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12635_ _05370_ _05374_ _05391_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__nand3_4
XFILLER_70_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15354_ _07968_ _08039_ vssd1 vssd1 vccd1 vccd1 _08040_ sky130_fd_sc_hd__xnor2_1
X_18142_ _04834_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__buf_4
XFILLER_184_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12566_ _05209_ _05322_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__nor2_4
XFILLER_196_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11517_ _04298_ _04299_ _03612_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__mux2_1
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14305_ _06992_ vssd1 vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__buf_4
XFILLER_184_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15285_ _07879_ _07884_ _07970_ vssd1 vssd1 vccd1 vccd1 _07971_ sky130_fd_sc_hd__a21bo_1
X_18073_ _02240_ vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12497_ _05158_ _05253_ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__or2_1
XFILLER_89_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19001__179 clknet_1_1__leaf__02731_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__inv_2
XFILLER_176_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17024_ _09606_ _09607_ vssd1 vssd1 vccd1 vccd1 _09629_ sky130_fd_sc_hd__or2_1
XFILLER_172_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14236_ _06922_ _06923_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__and2_1
X_11448_ _04231_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__inv_2
XFILLER_160_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14167_ _06854_ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__buf_6
XFILLER_98_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11379_ _04161_ _04162_ _03677_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__mux2_1
XFILLER_153_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13118_ _05873_ _05874_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__and2_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14098_ _05003_ vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__inv_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ _02162_ vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__clkbuf_1
X_13049_ _05484_ _05526_ _05805_ _05473_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__o22a_1
XFILLER_112_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17857_ rbzero.spi_registers.spi_counter\[4\] _01659_ rbzero.spi_registers.spi_counter\[6\]
+ rbzero.spi_registers.spi_counter\[5\] vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__a211oi_1
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16808_ _08485_ _09414_ _09415_ vssd1 vssd1 vccd1 vccd1 _09416_ sky130_fd_sc_hd__and3_2
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17788_ _01985_ rbzero.debug_overlay.vplaneX\[-2\] vssd1 vssd1 vccd1 vccd1 _02054_
+ sky130_fd_sc_hd__or2_1
XFILLER_81_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19527_ clknet_leaf_39_i_clk _00015_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[1\]
+ sky130_fd_sc_hd__dfxtp_4
X_16739_ _09345_ _09346_ vssd1 vssd1 vccd1 vccd1 _09347_ sky130_fd_sc_hd__xor2_1
XFILLER_35_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19458_ clknet_leaf_64_i_clk _00404_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19389_ _02860_ _02863_ _02864_ vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__and3_1
XFILLER_33_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20302_ net362 _01233_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20233_ net293 _01164_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18917__103 clknet_1_0__leaf__02723_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__inv_2
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09975_ _03041_ vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__clkbuf_1
X_20164_ net224 _01095_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20095_ clknet_leaf_90_i_clk _01026_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10750_ rbzero.color_sky\[0\] rbzero.color_floor\[0\] _03535_ vssd1 vssd1 vccd1 vccd1
+ _03536_ sky130_fd_sc_hd__mux2_1
X_18963__145 clknet_1_1__leaf__02727_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__inv_2
XFILLER_77_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10681_ gpout0.hpos\[3\] gpout0.hpos\[4\] gpout0.hpos\[5\] vssd1 vssd1 vccd1 vccd1
+ _03476_ sky130_fd_sc_hd__and3_1
XFILLER_198_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12420_ _05077_ _05150_ _05176_ _05152_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__a31o_1
XFILLER_138_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12351_ rbzero.wall_tracer.rcp_sel\[2\] _04898_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__nand2_1
XFILLER_181_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11302_ rbzero.debug_overlay.facingY\[-7\] _04083_ _04084_ rbzero.debug_overlay.facingY\[-6\]
+ _04086_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__a221o_1
XFILLER_193_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15070_ _07756_ _07199_ _07757_ _07185_ vssd1 vssd1 vccd1 vccd1 _07758_ sky130_fd_sc_hd__o22ai_1
XFILLER_14_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12282_ rbzero.debug_overlay.facingX\[-6\] rbzero.wall_tracer.rayAddendX\[2\] vssd1
+ vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__nor2_1
XFILLER_181_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14021_ _06664_ _06735_ vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__nand2_1
X_11233_ _04007_ _04010_ _04013_ _04017_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__or4_1
XFILLER_134_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11164_ rbzero.tex_r1\[39\] _03733_ _03948_ _03666_ vssd1 vssd1 vccd1 vccd1 _03949_
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10115_ rbzero.tex_g1\[9\] rbzero.tex_g1\[10\] _03106_ vssd1 vssd1 vccd1 vccd1 _03115_
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18760_ _02288_ _02632_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__and2_1
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11095_ rbzero.map_overlay.i_otherx\[0\] vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__inv_2
X_15972_ rbzero.wall_tracer.trackDistX\[-1\] rbzero.wall_tracer.stepDistX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _08587_ sky130_fd_sc_hd__nor2_1
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17711_ _01976_ _01982_ _03339_ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10046_ rbzero.tex_g1\[42\] rbzero.tex_g1\[43\] _03073_ vssd1 vssd1 vccd1 vccd1 _03079_
+ sky130_fd_sc_hd__mux2_1
X_14923_ _07574_ _07609_ vssd1 vssd1 vccd1 vccd1 _07611_ sky130_fd_sc_hd__xor2_1
X_18691_ rbzero.debug_overlay.playerY\[-9\] vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__inv_2
XFILLER_76_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17642_ rbzero.debug_overlay.vplaneX\[-6\] rbzero.wall_tracer.rayAddendX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__or2_1
X_14854_ _07536_ _07538_ vssd1 vssd1 vccd1 vccd1 _07542_ sky130_fd_sc_hd__or2_1
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13805_ _06330_ _06331_ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__or2_1
XFILLER_95_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17573_ _01784_ rbzero.debug_overlay.vplaneY\[-1\] vssd1 vssd1 vccd1 vccd1 _01860_
+ sky130_fd_sc_hd__and2_1
XFILLER_90_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11997_ _04750_ _04314_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__nand2_1
XFILLER_51_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14785_ _07374_ _07424_ vssd1 vssd1 vccd1 vccd1 _07473_ sky130_fd_sc_hd__or2_1
X_19312_ rbzero.traced_texa\[-2\] rbzero.texV\[-2\] vssd1 vssd1 vccd1 vccd1 _02800_
+ sky130_fd_sc_hd__or2_1
X_16524_ _06858_ _07012_ _07766_ _09133_ vssd1 vssd1 vccd1 vccd1 _09134_ sky130_fd_sc_hd__or4_1
XFILLER_1_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10948_ rbzero.tex_r0\[42\] _03733_ _03612_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__a21o_1
X_19081__251 clknet_1_0__leaf__02739_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__inv_2
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13736_ _06491_ _06486_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__and2b_1
XFILLER_189_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16455_ _09005_ _09065_ vssd1 vssd1 vccd1 vccd1 _09066_ sky130_fd_sc_hd__xnor2_1
X_10879_ rbzero.tex_r0\[15\] rbzero.tex_r0\[14\] _03664_ vssd1 vssd1 vccd1 vccd1 _03665_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13667_ _06398_ _06422_ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__and2b_1
XFILLER_188_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15406_ _08074_ _08090_ vssd1 vssd1 vccd1 vccd1 _08091_ sky130_fd_sc_hd__xor2_1
X_12618_ _05300_ _05308_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__and2_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16386_ _08861_ _08873_ _08871_ vssd1 vssd1 vccd1 vccd1 _08997_ sky130_fd_sc_hd__a21oi_1
X_13598_ _06307_ _06324_ vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__xnor2_1
XFILLER_185_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18125_ rbzero.spi_registers.new_other\[0\] _02264_ _02272_ _02266_ vssd1 vssd1 vccd1
+ vccd1 _00755_ sky130_fd_sc_hd__o211a_1
XFILLER_200_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15337_ _08012_ _08022_ vssd1 vssd1 vccd1 vccd1 _08023_ sky130_fd_sc_hd__xnor2_1
X_12549_ _05286_ _05290_ _05293_ _05296_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__or4b_2
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _03117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18056_ rbzero.spi_registers.spi_buffer\[4\] rbzero.spi_registers.spi_buffer\[3\]
+ _02227_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__mux2_1
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15268_ _07842_ _07785_ vssd1 vssd1 vccd1 vccd1 _07954_ sky130_fd_sc_hd__and2b_1
XFILLER_32_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17007_ _09611_ _09612_ vssd1 vssd1 vccd1 vccd1 _09613_ sky130_fd_sc_hd__nor2_1
XFILLER_132_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14219_ rbzero.wall_tracer.stepDistX\[-3\] vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__inv_2
X_15199_ _07876_ _07885_ vssd1 vssd1 vccd1 vccd1 _07886_ sky130_fd_sc_hd__xnor2_2
XFILLER_113_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09760_ rbzero.tex_r1\[48\] rbzero.tex_r1\[49\] _02921_ vssd1 vssd1 vccd1 vccd1 _02927_
+ sky130_fd_sc_hd__mux2_1
XFILLER_140_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17909_ rbzero.pov.spi_buffer\[9\] rbzero.pov.ready_buffer\[9\] _02153_ vssd1 vssd1
+ vccd1 vccd1 _02154_ sky130_fd_sc_hd__mux2_1
XFILLER_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18889_ _03902_ _02260_ _02713_ _02285_ vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__o211a_1
XFILLER_187_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19164__326 clknet_1_1__leaf__02747_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__inv_2
XFILLER_39_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20216_ net276 _01147_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20147_ clknet_leaf_13_i_clk _01078_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[5\] sky130_fd_sc_hd__dfxtp_4
XFILLER_104_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09958_ _03032_ vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20078_ clknet_leaf_7_i_clk _01009_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_09889_ _02996_ vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__clkbuf_1
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11920_ _03852_ _04672_ _04670_ _04694_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__a211o_1
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ net10 net9 vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__and2_1
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ rbzero.texV\[6\] _03586_ _03587_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__nand3_1
XFILLER_72_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _06866_ _07257_ vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__nor2_1
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11782_ net18 net19 vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__nand2_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13521_ _06228_ _06277_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__nor2_1
X_10733_ gpout0.vpos\[5\] gpout0.vpos\[4\] vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__or2_2
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16240_ _07984_ _07960_ _08070_ _07865_ vssd1 vssd1 vccd1 vccd1 _08852_ sky130_fd_sc_hd__o22a_1
X_13452_ _06205_ _06207_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__and2_1
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10664_ _02902_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__clkbuf_4
XFILLER_201_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12403_ rbzero.wall_tracer.visualWallDist\[6\] _03479_ vssd1 vssd1 vccd1 vccd1 _05160_
+ sky130_fd_sc_hd__nor2_1
XFILLER_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16171_ _08668_ _08765_ _08782_ vssd1 vssd1 vccd1 vccd1 _08784_ sky130_fd_sc_hd__nand3_1
XFILLER_127_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13383_ _06079_ _06139_ vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__xnor2_1
X_10595_ _03390_ _03358_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__nand2_1
XFILLER_103_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12334_ _05090_ _05083_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__xor2_2
X_15122_ _07808_ _07809_ vssd1 vssd1 vccd1 vccd1 _07810_ sky130_fd_sc_hd__nand2_1
XFILLER_193_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19930_ net159 _00861_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[10\] sky130_fd_sc_hd__dfxtp_1
X_15053_ _07728_ _07740_ vssd1 vssd1 vccd1 vccd1 _07741_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12265_ rbzero.wall_tracer.mapY\[9\] _04923_ _05019_ vssd1 vssd1 vccd1 vccd1 _05023_
+ sky130_fd_sc_hd__o21a_1
XFILLER_147_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14004_ _06747_ vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__clkbuf_1
X_11216_ rbzero.row_render.texu\[4\] _03688_ _03996_ vssd1 vssd1 vccd1 vccd1 _04001_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19861_ clknet_leaf_22_i_clk _00792_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12196_ rbzero.wall_tracer.trackDistY\[6\] vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__inv_2
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 o_hsync sky130_fd_sc_hd__buf_2
Xoutput71 net123 vssd1 vssd1 vccd1 vccd1 o_tex_sclk sky130_fd_sc_hd__clkbuf_1
X_18812_ rbzero.pov.ready_buffer\[32\] _02666_ _02667_ _02651_ vssd1 vssd1 vccd1 vccd1
+ _01047_ sky130_fd_sc_hd__a211o_1
X_11147_ rbzero.tex_r1\[61\] _03919_ _03926_ _03673_ vssd1 vssd1 vccd1 vccd1 _03932_
+ sky130_fd_sc_hd__a31o_1
XFILLER_122_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19792_ clknet_leaf_16_i_clk _00723_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18743_ _03337_ _02618_ _02622_ vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__or3_1
XFILLER_49_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11078_ rbzero.map_overlay.i_mapdx\[5\] _03421_ _03420_ vssd1 vssd1 vccd1 vccd1 _03864_
+ sky130_fd_sc_hd__o21a_1
X_15955_ _08563_ _08565_ _08564_ vssd1 vssd1 vccd1 vccd1 _08572_ sky130_fd_sc_hd__a21boi_1
XFILLER_95_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10029_ _03069_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__clkbuf_1
X_14906_ _07588_ _07593_ vssd1 vssd1 vccd1 vccd1 _07594_ sky130_fd_sc_hd__xor2_1
X_18674_ rbzero.debug_overlay.playerX\[2\] _02543_ _02569_ _02356_ vssd1 vssd1 vccd1
+ vccd1 _01007_ sky130_fd_sc_hd__o211a_1
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15886_ _07642_ _07691_ _08510_ vssd1 vssd1 vccd1 vccd1 _08511_ sky130_fd_sc_hd__o21a_1
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17625_ _04940_ _01904_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__xnor2_1
X_14837_ _07480_ _07524_ vssd1 vssd1 vccd1 vccd1 _07525_ sky130_fd_sc_hd__nor2_1
XFILLER_52_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17556_ _01827_ _01833_ _01842_ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__a21o_1
XFILLER_51_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14768_ _07429_ _07455_ vssd1 vssd1 vccd1 vccd1 _07456_ sky130_fd_sc_hd__xnor2_1
XFILLER_147_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16507_ _09115_ _09116_ vssd1 vssd1 vccd1 vccd1 _09117_ sky130_fd_sc_hd__xor2_1
XFILLER_149_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13719_ _06467_ _06466_ _06446_ vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17487_ _01762_ _01779_ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__xnor2_1
X_14699_ _07347_ _07384_ _07386_ _07344_ vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19007__185 clknet_1_0__leaf__02731_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__inv_2
XFILLER_176_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16438_ _09047_ _08803_ _09048_ vssd1 vssd1 vccd1 vccd1 _09049_ sky130_fd_sc_hd__or3b_1
XFILLER_176_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16369_ _08849_ _08853_ _08851_ vssd1 vssd1 vccd1 vccd1 _08980_ sky130_fd_sc_hd__a21oi_1
XFILLER_117_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18108_ _03852_ _02258_ _02260_ vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__and3_4
XFILLER_173_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18039_ _02221_ vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18992__171 clknet_1_0__leaf__02730_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__inv_2
XFILLER_160_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20001_ clknet_leaf_93_i_clk _00932_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_09812_ _02909_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__clkbuf_4
XFILLER_98_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09743_ rbzero.tex_r1\[56\] rbzero.tex_r1\[57\] _02910_ vssd1 vssd1 vccd1 vccd1 _02918_
+ sky130_fd_sc_hd__mux2_1
XFILLER_100_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19088__257 clknet_1_1__leaf__02740_ vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__inv_2
XFILLER_100_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10380_ _02908_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__clkbuf_4
XFILLER_109_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12050_ net36 net37 net38 _04822_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__or4_2
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11001_ rbzero.row_render.size\[3\] _03462_ _03463_ rbzero.row_render.size\[4\] _03786_
+ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__o221a_1
XFILLER_104_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19147__310 clknet_1_1__leaf__02746_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__inv_2
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15740_ _08421_ _08422_ vssd1 vssd1 vccd1 vccd1 _08423_ sky130_fd_sc_hd__nor2_1
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _05703_ _05708_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__xor2_1
XFILLER_92_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11903_ net22 _04670_ net24 vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__a21o_1
X_15671_ _08352_ _08353_ vssd1 vssd1 vccd1 vccd1 _08354_ sky130_fd_sc_hd__nand2_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _05633_ _05639_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ rbzero.debug_overlay.vplaneY\[-7\] rbzero.wall_tracer.rayAddendY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__nand2_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _07097_ _07100_ _07303_ vssd1 vssd1 vccd1 vccd1 _07310_ sky130_fd_sc_hd__or3_1
XFILLER_27_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _04571_ _04579_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__nand2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17341_ _01661_ vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__buf_2
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14553_ _07239_ _07240_ vssd1 vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__and2_1
X_11765_ gpout0.hpos\[0\] _03527_ _03526_ _04020_ net3 net4 vssd1 vssd1 vccd1 vccd1
+ _04543_ sky130_fd_sc_hd__mux4_1
XFILLER_198_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _06121_ _06035_ _06123_ vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__o21ai_1
X_10716_ _02900_ gpout0.hpos\[8\] gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 _03504_
+ sky130_fd_sc_hd__o21a_1
XFILLER_41_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17272_ rbzero.wall_tracer.trackDistY\[2\] rbzero.wall_tracer.stepDistY\[2\] vssd1
+ vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__nand2_1
XFILLER_201_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11696_ _04020_ _03464_ _03528_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__or3_1
X_14484_ _03492_ rbzero.wall_tracer.stepDistY\[4\] _04949_ vssd1 vssd1 vccd1 vccd1
+ _07172_ sky130_fd_sc_hd__a21oi_1
XFILLER_201_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16223_ rbzero.wall_tracer.trackDistX\[1\] rbzero.wall_tracer.stepDistX\[1\] vssd1
+ vssd1 vccd1 vccd1 _08836_ sky130_fd_sc_hd__nand2_1
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13435_ _06140_ _06191_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__nor2_1
X_10647_ rbzero.map_overlay.i_otherx\[1\] _03362_ rbzero.map_rom.i_col\[4\] _03441_
+ _03442_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__a221o_1
XFILLER_158_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16154_ _08000_ vssd1 vssd1 vccd1 vccd1 _08767_ sky130_fd_sc_hd__inv_2
X_19193__352 clknet_1_1__leaf__02750_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__inv_2
XFILLER_154_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13366_ _06002_ _06034_ _06054_ _06122_ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__a211o_1
XFILLER_127_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10578_ _03358_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__inv_2
X_15105_ _07782_ _07792_ vssd1 vssd1 vccd1 vccd1 _07793_ sky130_fd_sc_hd__nand2_1
XFILLER_177_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12317_ _05028_ _05058_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__nand2_1
XFILLER_177_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16085_ _08697_ _08698_ vssd1 vssd1 vccd1 vccd1 _08699_ sky130_fd_sc_hd__nor2_1
X_13297_ _06039_ _06033_ _06051_ _06053_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__a211oi_4
XFILLER_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15036_ _07125_ _07705_ _07723_ vssd1 vssd1 vccd1 vccd1 _07724_ sky130_fd_sc_hd__a21o_1
X_19913_ clknet_leaf_0_i_clk _00844_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12248_ _04945_ _05007_ _05008_ _05009_ rbzero.wall_tracer.mapY\[6\] vssd1 vssd1
+ vccd1 vccd1 _00401_ sky130_fd_sc_hd__a32o_1
XFILLER_130_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19844_ clknet_leaf_14_i_clk _00775_ vssd1 vssd1 vccd1 vccd1 rbzero.mapdyw\[0\] sky130_fd_sc_hd__dfxtp_1
X_12179_ _03375_ _04929_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__nand2_1
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19775_ clknet_leaf_5_i_clk _00706_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_16987_ _09577_ _09591_ vssd1 vssd1 vccd1 vccd1 _09593_ sky130_fd_sc_hd__or2_1
XFILLER_96_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18726_ rbzero.pov.ready_buffer\[53\] _02607_ _02540_ _02608_ _02581_ vssd1 vssd1
+ vccd1 vccd1 _02609_ sky130_fd_sc_hd__a221o_1
X_15938_ _08547_ _08549_ _08548_ vssd1 vssd1 vccd1 vccd1 _08557_ sky130_fd_sc_hd__a21boi_1
XFILLER_64_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18398__41 clknet_1_1__leaf__02435_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__inv_2
X_18657_ _02534_ _02555_ _02556_ _02356_ vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__o211a_1
X_15869_ _08493_ _08496_ vssd1 vssd1 vccd1 vccd1 _08497_ sky130_fd_sc_hd__xor2_1
XFILLER_149_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17608_ _01786_ _01888_ _01891_ _03484_ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18588_ _02513_ vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17539_ _01784_ rbzero.wall_tracer.rayAddendY\[5\] vssd1 vssd1 vccd1 vccd1 _01828_
+ sky130_fd_sc_hd__or2_1
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19209_ clknet_1_0__leaf__02743_ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__buf_1
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20481_ clknet_leaf_63_i_clk _01412_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09726_ _02899_ _02905_ _02907_ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__and3_2
XFILLER_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11550_ rbzero.tex_b0\[33\] rbzero.tex_b0\[32\] _03709_ vssd1 vssd1 vccd1 vccd1 _04332_
+ sky130_fd_sc_hd__mux2_1
XFILLER_129_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10501_ _03317_ vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11481_ _03661_ _04261_ _04262_ _04263_ _04198_ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__o221a_1
X_18999__177 clknet_1_1__leaf__02731_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__inv_2
XFILLER_109_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13220_ _05974_ _05976_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__xor2_2
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10432_ _03281_ vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13151_ _05857_ _05890_ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__nand2_1
XFILLER_163_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10363_ _03245_ vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12102_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] _04858_
+ _04862_ _04863_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__a221o_1
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13082_ _05489_ _05838_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__and2_1
X_10294_ rbzero.tex_b1\[52\] rbzero.tex_b1\[53\] _03199_ vssd1 vssd1 vccd1 vccd1 _03209_
+ sky130_fd_sc_hd__mux2_1
XFILLER_105_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16910_ _09515_ _09516_ vssd1 vssd1 vccd1 vccd1 _09517_ sky130_fd_sc_hd__and2b_1
X_12033_ _04797_ _04803_ _04805_ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__a21o_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17890_ rbzero.pov.spi_buffer\[0\] rbzero.pov.ready_buffer\[0\] _02143_ vssd1 vssd1
+ vccd1 vccd1 _02144_ sky130_fd_sc_hd__mux2_1
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16841_ _09446_ _09447_ vssd1 vssd1 vccd1 vccd1 _09448_ sky130_fd_sc_hd__nand2_1
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19560_ clknet_leaf_36_i_clk _00491_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.side
+ sky130_fd_sc_hd__dfxtp_4
X_16772_ _07992_ _09046_ vssd1 vssd1 vccd1 vccd1 _09380_ sky130_fd_sc_hd__nor2_1
XFILLER_59_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13984_ _05315_ _06728_ _06729_ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18511_ rbzero.pov.spi_buffer\[25\] rbzero.pov.spi_buffer\[26\] _02466_ vssd1 vssd1
+ vccd1 vccd1 _02473_ sky130_fd_sc_hd__mux2_1
X_15723_ _08403_ _08405_ vssd1 vssd1 vccd1 vccd1 _08406_ sky130_fd_sc_hd__xor2_2
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12935_ _05654_ _05690_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19491_ clknet_leaf_38_i_clk _00437_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15654_ _08097_ _08224_ vssd1 vssd1 vccd1 vccd1 _08337_ sky130_fd_sc_hd__nand2_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _05619_ _05580_ _05622_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__a21oi_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _07219_ _07226_ vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__xnor2_1
X_18373_ _02426_ _02415_ _02427_ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__and3b_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ net20 _04585_ _04592_ _04593_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__and4_1
XFILLER_15_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _04832_ _08267_ _08268_ _07162_ vssd1 vssd1 vccd1 vccd1 _08269_ sky130_fd_sc_hd__a31o_1
X_12797_ _05547_ _05553_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ rbzero.wall_tracer.trackDistY\[9\] rbzero.wall_tracer.stepDistY\[9\] vssd1
+ vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__or2_1
XFILLER_187_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14536_ _07078_ _06933_ _07221_ _07223_ vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__or4bb_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _04506_ _04511_ _04524_ _04525_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__a22o_2
XFILLER_109_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17255_ _01584_ _01585_ _01586_ vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__o21a_1
X_14467_ _07148_ _07154_ vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__or2_1
XFILLER_175_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11679_ rbzero.tex_b1\[7\] rbzero.tex_b1\[6\] _03699_ vssd1 vssd1 vccd1 vccd1 _04460_
+ sky130_fd_sc_hd__mux2_1
XFILLER_146_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16206_ _08660_ _08696_ _08818_ vssd1 vssd1 vccd1 vccd1 _08819_ sky130_fd_sc_hd__a21oi_2
X_13418_ _06168_ _06170_ _06174_ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__a21oi_1
X_17186_ rbzero.wall_tracer.trackDistY\[-11\] _01523_ _01528_ _08511_ vssd1 vssd1
+ vccd1 vccd1 _00560_ sky130_fd_sc_hd__o22a_1
X_14398_ _07083_ _07085_ _07082_ vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__a21bo_1
XFILLER_143_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16137_ _08640_ _08642_ _08748_ vssd1 vssd1 vccd1 vccd1 _08750_ sky130_fd_sc_hd__nand3_1
XFILLER_143_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13349_ _05616_ _06056_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__and2_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19119__286 clknet_1_1__leaf__02742_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__inv_2
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16068_ _07195_ _04950_ _07185_ _08399_ vssd1 vssd1 vccd1 vccd1 _08682_ sky130_fd_sc_hd__or4_2
XFILLER_64_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15019_ _06857_ _06979_ vssd1 vssd1 vccd1 vccd1 _07707_ sky130_fd_sc_hd__nor2_1
XFILLER_130_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19827_ clknet_leaf_13_i_clk _00758_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19758_ clknet_leaf_88_i_clk _00689_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18709_ _02596_ _06943_ _02539_ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__mux2_1
X_19689_ clknet_leaf_5_i_clk _00620_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.d6 sky130_fd_sc_hd__dfxtp_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20464_ net144 _01395_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20395_ net455 _01326_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10981_ _03620_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__buf_2
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12720_ _05210_ _05430_ _05431_ _05476_ _05432_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__a32o_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12651_ _05329_ _05405_ _05407_ _05269_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__a211o_1
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11602_ _03688_ _04357_ _04365_ _04383_ _03719_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__a311o_1
XFILLER_70_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12582_ _05336_ _05337_ _05338_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__a21oi_1
X_15370_ _08054_ _08055_ vssd1 vssd1 vccd1 vccd1 _08056_ sky130_fd_sc_hd__nand2_1
X_18392__36 clknet_1_1__leaf__02434_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__inv_2
XFILLER_184_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14321_ _06996_ _07008_ vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__or2b_1
X_11533_ rbzero.color_sky\[4\] rbzero.color_floor\[4\] _03535_ vssd1 vssd1 vccd1 vccd1
+ _04315_ sky130_fd_sc_hd__mux2_1
XFILLER_183_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17040_ _09643_ _09644_ vssd1 vssd1 vccd1 vccd1 _09645_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11464_ _03649_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__buf_6
X_14252_ _06939_ vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__clkbuf_4
XFILLER_137_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10415_ _03272_ vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__clkbuf_1
X_13203_ _05469_ _05918_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__or2_1
XFILLER_183_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11395_ _03669_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__buf_4
X_14183_ _04840_ rbzero.wall_tracer.stepDistX\[-10\] _06867_ _06870_ vssd1 vssd1 vccd1
+ vccd1 _06871_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_174_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10346_ _03236_ vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__clkbuf_1
X_13134_ _05857_ _05890_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__xnor2_1
XFILLER_152_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17942_ rbzero.pov.spi_buffer\[25\] rbzero.pov.ready_buffer\[25\] _02164_ vssd1 vssd1
+ vccd1 vccd1 _02171_ sky130_fd_sc_hd__mux2_1
X_13065_ _05818_ _05809_ _05817_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__and3_1
X_10277_ _03200_ vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__clkbuf_1
X_12016_ net38 _04788_ net34 net35 vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__and4b_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17873_ rbzero.spi_registers.spi_counter\[2\] rbzero.spi_registers.spi_counter\[1\]
+ rbzero.spi_registers.spi_counter\[0\] rbzero.spi_registers.spi_counter\[3\] vssd1
+ vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__a31o_1
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16824_ _09374_ _09355_ vssd1 vssd1 vccd1 vccd1 _09431_ sky130_fd_sc_hd__or2b_1
X_19612_ clknet_leaf_53_i_clk _00543_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19543_ clknet_leaf_67_i_clk _00474_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.side
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_81_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16755_ _09016_ _09035_ _09036_ _09014_ vssd1 vssd1 vccd1 vccd1 _09363_ sky130_fd_sc_hd__o22ai_1
XFILLER_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13967_ _06665_ _06683_ _06699_ _06714_ _05380_ _05310_ vssd1 vssd1 vccd1 vccd1 _06715_
+ sky130_fd_sc_hd__mux4_2
XFILLER_98_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15706_ _07661_ _08260_ vssd1 vssd1 vccd1 vccd1 _08389_ sky130_fd_sc_hd__nor2_1
XFILLER_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12918_ _05665_ _05674_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__xor2_1
XFILLER_62_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19474_ clknet_leaf_50_i_clk _00420_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16686_ _09293_ _09294_ vssd1 vssd1 vccd1 vccd1 _09295_ sky130_fd_sc_hd__nor2_1
XFILLER_62_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13898_ _06603_ _06625_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__nor2_1
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15637_ _07672_ _08314_ _08315_ _08319_ vssd1 vssd1 vccd1 vccd1 _08320_ sky130_fd_sc_hd__o31a_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _05355_ _05496_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__nor2_2
XFILLER_61_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19125__290 clknet_1_0__leaf__02744_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__inv_2
X_18356_ rbzero.pov.ss_buffer\[1\] _02981_ vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__nor2_2
X_15568_ _07137_ vssd1 vssd1 vccd1 vccd1 _08252_ sky130_fd_sc_hd__buf_2
XFILLER_159_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17307_ _01534_ _01631_ _01632_ _01526_ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__a31o_1
X_14519_ _07189_ _07205_ vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__nand2_1
XFILLER_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18287_ rbzero.spi_registers.spi_buffer\[5\] rbzero.spi_registers.new_floor\[5\]
+ _02370_ vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__mux2_1
X_15499_ _08170_ _08171_ vssd1 vssd1 vccd1 vccd1 _08183_ sky130_fd_sc_hd__nor2_1
XFILLER_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17238_ rbzero.wall_tracer.trackDistY\[-3\] rbzero.wall_tracer.stepDistY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__and2_1
XFILLER_70_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17169_ _01457_ _01512_ _08509_ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__a21oi_1
XFILLER_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20180_ net240 _01111_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09991_ _03049_ vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20516_ clknet_leaf_77_i_clk _01447_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20447_ net507 _01378_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[38\] sky130_fd_sc_hd__dfxtp_1
X_10200_ rbzero.tex_g0\[34\] rbzero.tex_g0\[33\] _03155_ vssd1 vssd1 vccd1 vccd1 _03160_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11180_ rbzero.tex_r1\[1\] _03660_ _03768_ _03670_ vssd1 vssd1 vccd1 vccd1 _03965_
+ sky130_fd_sc_hd__a31o_1
XFILLER_107_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20378_ net438 _01309_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10131_ _03123_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10062_ _03087_ vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14870_ _07553_ _07557_ vssd1 vssd1 vccd1 vccd1 _07558_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13821_ _06196_ _06576_ _06577_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__nor3b_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16540_ _09042_ _09132_ _09149_ vssd1 vssd1 vccd1 vccd1 _09150_ sky130_fd_sc_hd__a21o_1
X_13752_ _06477_ _06508_ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__and2_1
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10964_ rbzero.tex_r0\[61\] rbzero.tex_r0\[60\] _03663_ vssd1 vssd1 vccd1 vccd1 _03750_
+ sky130_fd_sc_hd__mux2_1
X_12703_ _05367_ _05405_ _05435_ _05270_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__o211ai_1
X_16471_ rbzero.wall_tracer.trackDistX\[3\] rbzero.wall_tracer.stepDistX\[3\] vssd1
+ vssd1 vccd1 vccd1 _09082_ sky130_fd_sc_hd__nand2_1
X_13683_ _05862_ _06035_ _06439_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__or3b_1
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10895_ _03589_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__inv_2
X_18210_ _02327_ vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__clkbuf_1
X_15422_ _07097_ vssd1 vssd1 vccd1 vccd1 _08107_ sky130_fd_sc_hd__clkbuf_4
XFILLER_31_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12634_ _05376_ _05381_ _05389_ _05390_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__a211o_1
XFILLER_93_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18940__124 clknet_1_0__leaf__02725_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__inv_2
XFILLER_54_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18141_ rbzero.spi_registers.got_new_vinf _02262_ rbzero.row_render.vinf vssd1 vssd1
+ vccd1 vccd1 _02284_ sky130_fd_sc_hd__a21o_1
XFILLER_141_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15353_ _08036_ _08038_ vssd1 vssd1 vccd1 vccd1 _08039_ sky130_fd_sc_hd__xor2_1
XFILLER_54_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12565_ _05321_ _05300_ _05278_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__a21boi_4
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14304_ _06984_ _06986_ _06991_ _04948_ vssd1 vssd1 vccd1 vccd1 _06992_ sky130_fd_sc_hd__a22o_1
X_11516_ rbzero.tex_g1\[41\] rbzero.tex_g1\[40\] _03727_ vssd1 vssd1 vccd1 vccd1 _04299_
+ sky130_fd_sc_hd__mux2_1
X_18072_ rbzero.spi_registers.spi_buffer\[12\] rbzero.spi_registers.spi_buffer\[11\]
+ _02226_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__mux2_1
X_15284_ _07885_ _07876_ vssd1 vssd1 vccd1 vccd1 _07970_ sky130_fd_sc_hd__or2b_1
XFILLER_102_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12496_ _05204_ _05206_ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__or2_1
XFILLER_184_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17023_ _09622_ _09628_ rbzero.wall_tracer.trackDistX\[8\] _08508_ vssd1 vssd1 vccd1
+ vccd1 _00557_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_176_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14235_ rbzero.debug_overlay.playerY\[-6\] _06877_ vssd1 vssd1 vccd1 vccd1 _06923_
+ sky130_fd_sc_hd__nand2_1
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11447_ _03896_ _03847_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__or2_1
X_11378_ rbzero.tex_g0\[27\] rbzero.tex_g0\[26\] _03709_ vssd1 vssd1 vccd1 vccd1 _04162_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14166_ rbzero.wall_tracer.state\[6\] rbzero.wall_tracer.state\[13\] vssd1 vssd1
+ vccd1 vccd1 _06854_ sky130_fd_sc_hd__nor2_2
XFILLER_140_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10329_ _03227_ vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__clkbuf_1
X_13117_ _05859_ _05860_ _05872_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__nand3_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ rbzero.wall_tracer.trackDistX\[10\] _04953_ rbzero.wall_tracer.trackDistY\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__o21a_1
XFILLER_140_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17925_ rbzero.pov.spi_buffer\[17\] rbzero.pov.ready_buffer\[17\] _02153_ vssd1 vssd1
+ vccd1 vccd1 _02162_ sky130_fd_sc_hd__mux2_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _05535_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__clkbuf_4
XFILLER_39_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17856_ _01659_ _02105_ _02106_ _02109_ _02116_ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__o311a_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16807_ _09410_ _09413_ vssd1 vssd1 vccd1 vccd1 _09415_ sky130_fd_sc_hd__or2_1
XFILLER_54_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17787_ _02050_ _02051_ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__or2_1
X_14999_ _07645_ _07685_ _07666_ _07650_ vssd1 vssd1 vccd1 vccd1 _07687_ sky130_fd_sc_hd__a211o_1
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16738_ _09227_ _09239_ _09237_ vssd1 vssd1 vccd1 vccd1 _09346_ sky130_fd_sc_hd__a21oi_1
X_19526_ clknet_leaf_67_i_clk _00013_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19457_ clknet_leaf_64_i_clk _00403_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16669_ _09268_ _09276_ vssd1 vssd1 vccd1 vccd1 _09278_ sky130_fd_sc_hd__or2_1
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19388_ rbzero.traced_texa\[10\] rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 _02864_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_194_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18339_ rbzero.spi_registers.new_vshift\[3\] rbzero.spi_registers.spi_buffer\[3\]
+ _02401_ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__mux2_1
XFILLER_147_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20301_ net361 _01232_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20232_ net292 _01163_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20163_ net223 _01094_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09974_ rbzero.tex_r0\[13\] rbzero.tex_r0\[12\] _03039_ vssd1 vssd1 vccd1 vccd1 _03041_
+ sky130_fd_sc_hd__mux2_1
XFILLER_157_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20094_ clknet_leaf_8_i_clk _01025_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_57_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_54_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_69_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19141__305 clknet_1_1__leaf__02745_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__inv_2
XFILLER_164_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10680_ _02901_ _03474_ _02902_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__or3_1
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12350_ _05040_ _05106_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__xnor2_4
X_11301_ rbzero.debug_overlay.facingY\[-5\] _04085_ _03900_ _03849_ vssd1 vssd1 vccd1
+ vccd1 _04086_ sky130_fd_sc_hd__a211o_1
XFILLER_154_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12281_ rbzero.debug_overlay.facingX\[-7\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__nor2_1
XFILLER_153_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11232_ _03902_ _03461_ _04016_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__a21oi_1
X_14020_ _05315_ _06723_ vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__nand2_1
XFILLER_101_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11163_ rbzero.tex_r1\[38\] _03767_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__or2_1
XFILLER_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10114_ _03114_ vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11094_ gpout0.vpos\[3\] rbzero.map_overlay.i_othery\[0\] vssd1 vssd1 vccd1 vccd1
+ _03880_ sky130_fd_sc_hd__or2_1
X_15971_ rbzero.wall_tracer.trackDistX\[-1\] rbzero.wall_tracer.stepDistX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _08586_ sky130_fd_sc_hd__and2_1
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17710_ _01979_ _01981_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10045_ _03078_ vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14922_ _07574_ _07609_ vssd1 vssd1 vccd1 vccd1 _07610_ sky130_fd_sc_hd__and2_1
X_18690_ _02581_ vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__buf_2
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17641_ _01916_ _01917_ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__and2b_1
XFILLER_64_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14853_ _07540_ vssd1 vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__clkbuf_2
XFILLER_36_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13804_ _06335_ _06431_ _06434_ _06560_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__a22o_1
X_17572_ _01785_ rbzero.debug_overlay.vplaneY\[-1\] vssd1 vssd1 vccd1 vccd1 _01859_
+ sky130_fd_sc_hd__nor2_1
X_14784_ _07365_ _07367_ vssd1 vssd1 vccd1 vccd1 _07472_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11996_ _04741_ _04758_ _04769_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__and3_2
XFILLER_1_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19311_ _02759_ _02798_ _02799_ _02762_ rbzero.texV\[-3\] vssd1 vssd1 vccd1 vccd1
+ _01414_ sky130_fd_sc_hd__a32o_1
X_16523_ _08130_ vssd1 vssd1 vccd1 vccd1 _09133_ sky130_fd_sc_hd__buf_2
XFILLER_44_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13735_ _06486_ _06491_ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__and2b_1
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10947_ _03732_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__clkbuf_4
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19242_ clknet_1_0__leaf__04486_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__buf_1
X_16454_ _09063_ _09064_ vssd1 vssd1 vccd1 vccd1 _09065_ sky130_fd_sc_hd__and2b_1
XFILLER_32_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13666_ _06398_ _06422_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__xnor2_1
X_10878_ _03663_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__buf_4
XFILLER_176_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15405_ _08087_ _08089_ vssd1 vssd1 vccd1 vccd1 _08090_ sky130_fd_sc_hd__xor2_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _05371_ _05372_ _05373_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__o21ai_2
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16385_ _08986_ _08995_ vssd1 vssd1 vccd1 vccd1 _08996_ sky130_fd_sc_hd__xnor2_1
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13597_ _06342_ _06351_ _06353_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__a21oi_2
XFILLER_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18124_ _03437_ _02263_ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__nand2_1
X_15336_ _07900_ _08019_ _08021_ vssd1 vssd1 vccd1 vccd1 _08022_ sky130_fd_sc_hd__a21oi_1
XFILLER_185_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12548_ _05234_ _05243_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__nor2_2
XFILLER_200_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18055_ _02231_ vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__clkbuf_1
X_15267_ _07951_ _07952_ vssd1 vssd1 vccd1 vccd1 _07953_ sky130_fd_sc_hd__nand2_1
XFILLER_172_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12479_ _03489_ _05107_ _05109_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__a21oi_2
XANTENNA_2 _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17006_ _09318_ _09513_ _09511_ vssd1 vssd1 vccd1 vccd1 _09612_ sky130_fd_sc_hd__a21oi_1
XFILLER_144_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14218_ _04947_ vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__buf_4
XFILLER_99_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15198_ _07879_ _07884_ vssd1 vssd1 vccd1 vccd1 _07885_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14149_ _03455_ _03389_ vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__or2b_1
XFILLER_113_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17908_ _02142_ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__clkbuf_4
XFILLER_39_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18888_ _02712_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__inv_2
XFILLER_94_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17839_ _01714_ _02099_ _02100_ _08458_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__o22a_1
XFILLER_55_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19509_ clknet_leaf_58_i_clk _00455_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20215_ net275 _01146_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20146_ clknet_leaf_13_i_clk _01077_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[4\] sky130_fd_sc_hd__dfxtp_1
X_09957_ rbzero.tex_r0\[21\] rbzero.tex_r0\[20\] _03028_ vssd1 vssd1 vccd1 vccd1 _03032_
+ sky130_fd_sc_hd__mux2_1
XFILLER_103_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20077_ clknet_leaf_86_i_clk _01008_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_09888_ rbzero.tex_r0\[54\] rbzero.tex_r0\[53\] _02995_ vssd1 vssd1 vccd1 vccd1 _02996_
+ sky130_fd_sc_hd__mux2_1
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ net9 net10 vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__and2b_1
XFILLER_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10801_ rbzero.traced_texVinit\[6\] rbzero.spi_registers.vshift\[3\] vssd1 vssd1
+ vccd1 vccd1 _03587_ sky130_fd_sc_hd__or2_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _04552_ _04393_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__nor2_1
XFILLER_199_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13520_ _06229_ _06272_ _06276_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__o21a_1
XFILLER_198_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10732_ gpout0.vpos\[2\] gpout0.vpos\[1\] gpout0.vpos\[0\] vssd1 vssd1 vccd1 vccd1
+ _03518_ sky130_fd_sc_hd__or3_2
XFILLER_198_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13451_ _06205_ _06207_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__nor2_1
XFILLER_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10663_ _03340_ _03458_ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__nor2_2
XFILLER_90_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12402_ _05077_ _05150_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__and2_1
XFILLER_185_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16170_ _08668_ _08765_ _08782_ vssd1 vssd1 vccd1 vccd1 _08783_ sky130_fd_sc_hd__a21o_1
XFILLER_166_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10594_ rbzero.map_rom.d6 vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__clkbuf_4
X_13382_ _06116_ _06138_ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__xor2_1
XFILLER_182_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15121_ rbzero.debug_overlay.playerY\[-6\] rbzero.debug_overlay.playerX\[-6\] _06851_
+ vssd1 vssd1 vccd1 vccd1 _07809_ sky130_fd_sc_hd__mux2_1
X_12333_ _05084_ _05052_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__nand2_1
XFILLER_193_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15052_ _07738_ _07739_ vssd1 vssd1 vccd1 vccd1 _07740_ sky130_fd_sc_hd__nand2_1
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12264_ _05007_ _05021_ _05022_ _05009_ rbzero.wall_tracer.mapY\[9\] vssd1 vssd1
+ vccd1 vccd1 _00404_ sky130_fd_sc_hd__a32o_1
XFILLER_123_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14003_ rbzero.wall_tracer.stepDistY\[2\] _06746_ _06718_ vssd1 vssd1 vccd1 vccd1
+ _06747_ sky130_fd_sc_hd__mux2_1
XFILLER_141_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11215_ rbzero.row_render.texu\[4\] _03687_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__or2_1
XFILLER_107_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12195_ rbzero.wall_tracer.trackDistY\[7\] vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__inv_2
X_19860_ clknet_leaf_23_i_clk _00791_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 o_reset sky130_fd_sc_hd__buf_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 o_vsync sky130_fd_sc_hd__buf_2
X_18811_ rbzero.debug_overlay.facingY\[10\] _02634_ vssd1 vssd1 vccd1 vccd1 _02667_
+ sky130_fd_sc_hd__and2_1
X_11146_ rbzero.tex_r1\[63\] _03925_ _03930_ _03917_ vssd1 vssd1 vccd1 vccd1 _03931_
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19791_ clknet_leaf_7_i_clk _00722_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_122_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18742_ rbzero.pov.ready_buffer\[56\] _02539_ _02620_ _02621_ _02587_ vssd1 vssd1
+ vccd1 vccd1 _02622_ sky130_fd_sc_hd__o221a_1
X_11077_ _03425_ _03523_ _03464_ rbzero.map_overlay.i_mapdx\[1\] _03862_ vssd1 vssd1
+ vccd1 vccd1 _03863_ sky130_fd_sc_hd__a221o_1
X_15954_ _08569_ _06907_ vssd1 vssd1 vccd1 vccd1 _08571_ sky130_fd_sc_hd__nor2_1
XFILLER_95_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10028_ rbzero.tex_g1\[50\] rbzero.tex_g1\[51\] _03061_ vssd1 vssd1 vccd1 vccd1 _03069_
+ sky130_fd_sc_hd__mux2_1
X_14905_ _07589_ _07592_ _07590_ vssd1 vssd1 vccd1 vccd1 _07593_ sky130_fd_sc_hd__o21a_1
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18673_ rbzero.pov.ready_buffer\[70\] _02413_ _02533_ _02568_ vssd1 vssd1 vccd1 vccd1
+ _02569_ sky130_fd_sc_hd__a211o_1
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15885_ _07642_ _07691_ _08509_ vssd1 vssd1 vccd1 vccd1 _08510_ sky130_fd_sc_hd__a21oi_1
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17624_ _04941_ _01903_ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__nand2_1
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14836_ _07497_ _07522_ _07523_ vssd1 vssd1 vccd1 vccd1 _07524_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ _01827_ _01833_ _01842_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__nand3_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14767_ _07430_ _07431_ vssd1 vssd1 vccd1 vccd1 _07455_ sky130_fd_sc_hd__and2b_1
X_11979_ _04503_ _04750_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__nor2_1
XFILLER_44_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16506_ _07993_ _08081_ vssd1 vssd1 vccd1 vccd1 _09116_ sky130_fd_sc_hd__nor2_1
XFILLER_177_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13718_ _06446_ _06467_ _06466_ vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__and3_1
XFILLER_147_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17486_ _01777_ _01778_ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__nor2_1
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14698_ rbzero.wall_tracer.visualWallDist\[-10\] _04839_ _06985_ _06905_ vssd1 vssd1
+ vccd1 vccd1 _07386_ sky130_fd_sc_hd__and4_1
XFILLER_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16437_ _07617_ _07646_ _08681_ vssd1 vssd1 vccd1 vccd1 _09048_ sky130_fd_sc_hd__or3_2
XFILLER_20_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13649_ _06388_ _06405_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__nor2_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16368_ _08975_ _08978_ vssd1 vssd1 vccd1 vccd1 _08979_ sky130_fd_sc_hd__xor2_1
XFILLER_145_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18107_ _03834_ _03506_ _02259_ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__and3_1
X_15319_ _07881_ _07994_ _08003_ vssd1 vssd1 vccd1 vccd1 _08005_ sky130_fd_sc_hd__nand3_1
XFILLER_9_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19087_ clknet_1_1__leaf__02732_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__buf_1
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16299_ _07581_ _07897_ vssd1 vssd1 vccd1 vccd1 _08911_ sky130_fd_sc_hd__nor2_1
X_18038_ rbzero.pov.spi_buffer\[71\] rbzero.pov.ready_buffer\[71\] _02142_ vssd1 vssd1
+ vccd1 vccd1 _02221_ sky130_fd_sc_hd__mux2_1
XFILLER_105_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19170__331 clknet_1_0__leaf__02748_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__inv_2
XFILLER_67_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20000_ clknet_leaf_93_i_clk _00931_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_09811_ _02953_ vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19989_ clknet_leaf_95_i_clk _00920_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09742_ _02917_ vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11000_ rbzero.row_render.size\[2\] _03783_ _03462_ rbzero.row_render.size\[3\] _03785_
+ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__a221o_1
XFILLER_81_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20129_ clknet_leaf_89_i_clk _01060_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_86_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ _05704_ _05707_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__nand2_1
XFILLER_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11902_ _04667_ _04671_ _04676_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__o21a_1
X_15670_ _08240_ _08324_ _08351_ vssd1 vssd1 vccd1 vccd1 _08353_ sky130_fd_sc_hd__nand3_1
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _05636_ _05638_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__and2_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _06971_ _06994_ _06967_ vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__a21bo_1
XFILLER_73_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ net20 _04563_ _04583_ _04609_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__a31o_2
XFILLER_27_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17340_ rbzero.spi_registers.spi_done _02907_ _01660_ vssd1 vssd1 vccd1 vccd1 _01661_
+ sky130_fd_sc_hd__and3_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _07223_ _07224_ _07238_ vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__nand3_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _03459_ _03469_ net3 vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__mux2_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13503_ _06171_ _06173_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__xnor2_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _03462_ _03502_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__nor2_1
XFILLER_92_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17271_ rbzero.wall_tracer.trackDistY\[1\] _01558_ _01601_ _08835_ vssd1 vssd1 vccd1
+ vccd1 _00572_ sky130_fd_sc_hd__o22a_1
XFILLER_186_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14483_ _04831_ _07169_ _07170_ _07162_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__a31o_1
X_11695_ _02899_ _04032_ _03528_ _04474_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__a31o_1
X_19010_ clknet_1_1__leaf__02732_ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__buf_1
XFILLER_158_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16222_ _08524_ _08834_ vssd1 vssd1 vccd1 vccd1 _08835_ sky130_fd_sc_hd__and2_1
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13434_ _06165_ _06190_ _06188_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__a21oi_1
XFILLER_186_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10646_ rbzero.map_overlay.i_otherx\[0\] _03395_ vssd1 vssd1 vccd1 vccd1 _03442_
+ sky130_fd_sc_hd__xor2_1
X_16153_ rbzero.wall_tracer.visualWallDist\[1\] _07256_ vssd1 vssd1 vccd1 vccd1 _08766_
+ sky130_fd_sc_hd__and2_1
XFILLER_154_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13365_ _05536_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__buf_2
XFILLER_158_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10577_ rbzero.map_rom.f4 vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__inv_2
X_15104_ _07790_ _07791_ vssd1 vssd1 vccd1 vccd1 _07792_ sky130_fd_sc_hd__and2_1
XFILLER_127_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12316_ _05029_ _05057_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__nand2_1
X_16084_ _08377_ _08414_ _08413_ vssd1 vssd1 vccd1 vccd1 _08698_ sky130_fd_sc_hd__a21oi_2
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13296_ _06004_ _06052_ _06032_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__a21boi_1
XFILLER_114_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15035_ _07712_ _07722_ vssd1 vssd1 vccd1 vccd1 _07723_ sky130_fd_sc_hd__xnor2_1
X_19912_ clknet_leaf_7_i_clk _00843_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready sky130_fd_sc_hd__dfxtp_1
X_12247_ _05006_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__clkbuf_4
XFILLER_111_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19843_ clknet_leaf_17_i_clk _00774_ vssd1 vssd1 vccd1 vccd1 rbzero.mapdxw\[1\] sky130_fd_sc_hd__dfxtp_1
X_12178_ _04936_ _04939_ _04937_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__a21o_1
XFILLER_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11129_ rbzero.color_floor\[1\] _03535_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__or2b_1
X_19774_ clknet_leaf_5_i_clk _00705_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_16986_ _09577_ _09591_ vssd1 vssd1 vccd1 vccd1 _09592_ sky130_fd_sc_hd__nand2_1
XFILLER_77_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18725_ rbzero.debug_overlay.playerY\[0\] _07026_ vssd1 vssd1 vccd1 vccd1 _02608_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_83_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15937_ rbzero.wall_tracer.trackDistX\[-5\] rbzero.wall_tracer.stepDistX\[-5\] vssd1
+ vssd1 vccd1 vccd1 _08556_ sky130_fd_sc_hd__and2_1
XFILLER_149_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18656_ _07022_ _02533_ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__nand2_1
X_15868_ _08467_ _08494_ _08495_ vssd1 vssd1 vccd1 vccd1 _08496_ sky130_fd_sc_hd__or3_1
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17607_ _01889_ _01890_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__xnor2_1
X_14819_ _07451_ _07505_ _07506_ vssd1 vssd1 vccd1 vccd1 _07507_ sky130_fd_sc_hd__a21oi_2
XFILLER_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18587_ rbzero.pov.spi_buffer\[61\] rbzero.pov.spi_buffer\[62\] _02510_ vssd1 vssd1
+ vccd1 vccd1 _02513_ sky130_fd_sc_hd__mux2_1
X_15799_ rbzero.row_render.texu\[2\] _08456_ _08453_ rbzero.wall_tracer.texu\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__a22o_1
X_17538_ _01784_ rbzero.wall_tracer.rayAddendY\[5\] vssd1 vssd1 vccd1 vccd1 _01827_
+ sky130_fd_sc_hd__nand2_1
XFILLER_33_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17469_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.debug_overlay.vplaneY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__nand2_1
XFILLER_193_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20480_ clknet_leaf_62_i_clk _01411_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09725_ _02906_ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__buf_6
XFILLER_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10500_ rbzero.tex_b0\[19\] rbzero.tex_b0\[18\] _03313_ vssd1 vssd1 vccd1 vccd1 _03317_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19177__337 clknet_1_1__leaf__02749_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__inv_2
X_11480_ rbzero.tex_g1\[9\] _03729_ _03730_ _03917_ vssd1 vssd1 vccd1 vccd1 _04263_
+ sky130_fd_sc_hd__a31o_1
XFILLER_149_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10431_ rbzero.tex_b0\[52\] rbzero.tex_b0\[51\] _03280_ vssd1 vssd1 vccd1 vccd1 _03281_
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13150_ _05894_ _05897_ _05899_ _05856_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__a2bb2o_1
X_10362_ rbzero.tex_b1\[20\] rbzero.tex_b1\[21\] _03243_ vssd1 vssd1 vccd1 vccd1 _03245_
+ sky130_fd_sc_hd__mux2_1
XFILLER_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12101_ rbzero.debug_overlay.facingY\[-7\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__and2_1
X_10293_ _03208_ vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__clkbuf_1
X_13081_ _05558_ _05806_ _05808_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__a21oi_1
XFILLER_151_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12032_ net36 net35 _04804_ net37 vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__a31o_1
XFILLER_104_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16840_ _09133_ _09231_ _09337_ vssd1 vssd1 vccd1 vccd1 _09447_ sky130_fd_sc_hd__o21bai_1
XFILLER_78_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16771_ _09377_ _09378_ vssd1 vssd1 vccd1 vccd1 _09379_ sky130_fd_sc_hd__and2_1
X_13983_ _05380_ _06714_ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__or2_1
X_15722_ _08145_ _08270_ _08404_ vssd1 vssd1 vccd1 vccd1 _08405_ sky130_fd_sc_hd__a21o_1
X_18510_ _02472_ vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__clkbuf_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12934_ _05526_ _05474_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__or2_1
XFILLER_74_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19490_ clknet_leaf_61_i_clk _00436_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15653_ _07856_ _08081_ _08208_ _08207_ vssd1 vssd1 vccd1 vccd1 _08336_ sky130_fd_sc_hd__o31ai_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ _05616_ _05620_ _05621_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__mux2_1
XFILLER_18_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _07231_ _07242_ vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__xnor2_1
XFILLER_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ rbzero.pov.spi_counter\[3\] rbzero.pov.spi_counter\[2\] _02417_ rbzero.pov.spi_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__a31o_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ net18 net17 net19 vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__a21o_1
XFILLER_57_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _06771_ _06776_ _07893_ _08266_ vssd1 vssd1 vccd1 vccd1 _08268_ sky130_fd_sc_hd__a31o_1
X_12796_ _05492_ _05548_ _05552_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__a21oi_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ rbzero.wall_tracer.trackDistY\[9\] rbzero.wall_tracer.stepDistY\[9\] vssd1
+ vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__nand2_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _07118_ _07222_ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__or2_1
XFILLER_30_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ net8 net7 vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__nor2_1
XFILLER_187_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17254_ _01584_ _01585_ _01586_ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__nor3_1
XFILLER_119_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14466_ _04949_ rbzero.wall_tracer.stepDistX\[2\] _07152_ _07153_ vssd1 vssd1 vccd1
+ vccd1 _07154_ sky130_fd_sc_hd__a22oi_4
X_11678_ rbzero.tex_b1\[5\] rbzero.tex_b1\[4\] _03699_ vssd1 vssd1 vccd1 vccd1 _04459_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16205_ _08693_ _08695_ vssd1 vssd1 vccd1 vccd1 _08818_ sky130_fd_sc_hd__nor2_1
XFILLER_30_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13417_ _06171_ _06173_ vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__and2_1
X_10629_ rbzero.map_overlay.i_mapdx\[0\] vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__inv_2
X_17185_ _08562_ _01524_ _01525_ _01527_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__a31o_1
X_14397_ _07084_ _06993_ vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__nor2_1
XFILLER_183_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16136_ _08640_ _08642_ _08748_ vssd1 vssd1 vccd1 vccd1 _08749_ sky130_fd_sc_hd__a21o_1
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13348_ _06087_ _06088_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__nand2_1
XFILLER_185_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16067_ _08396_ _08399_ vssd1 vssd1 vccd1 vccd1 _08681_ sky130_fd_sc_hd__or2_2
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13279_ _06001_ _05987_ _06035_ _05503_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__o22a_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15018_ _06875_ _07007_ vssd1 vssd1 vccd1 vccd1 _07706_ sky130_fd_sc_hd__nor2_1
XFILLER_64_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19826_ clknet_leaf_19_i_clk _00757_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19757_ clknet_leaf_88_i_clk _00688_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_56_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16969_ _09573_ _09574_ vssd1 vssd1 vccd1 vccd1 _09575_ sky130_fd_sc_hd__nor2_1
XFILLER_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18708_ rbzero.pov.ready_buffer\[48\] vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__inv_2
X_19688_ clknet_leaf_67_i_clk _00619_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18639_ _02534_ _02541_ _02544_ _02356_ vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__o211a_1
XFILLER_80_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20463_ net143 _01394_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20394_ net454 _01325_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10980_ _03537_ _03541_ _03647_ _03765_ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__a31o_1
XFILLER_74_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12650_ _05294_ _05313_ _05406_ _05304_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__o211a_1
XFILLER_31_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11601_ _03679_ _04369_ _04373_ _03684_ _04382_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__o311a_1
X_12581_ _05304_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__clkbuf_4
XFILLER_169_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14320_ _06997_ _07000_ _07007_ _06999_ vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__o31ai_2
XFILLER_12_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11532_ _04314_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkinv_2
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ _06938_ vssd1 vssd1 vccd1 vccd1 _06939_ sky130_fd_sc_hd__buf_2
XFILLER_183_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11463_ _04242_ _04245_ _03671_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__mux2_1
XFILLER_171_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13202_ _05957_ _05958_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__or2_1
X_10414_ rbzero.tex_b0\[60\] rbzero.tex_b0\[59\] _03269_ vssd1 vssd1 vccd1 vccd1 _03272_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14182_ _06853_ _06649_ _06869_ vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__o21ai_1
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11394_ _03739_ _04177_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__or2_1
XFILLER_178_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13133_ _05888_ _05889_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__and2_1
X_10345_ rbzero.tex_b1\[28\] rbzero.tex_b1\[29\] _03232_ vssd1 vssd1 vccd1 vccd1 _03236_
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13064_ _05728_ _05820_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__xor2_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17941_ _02170_ vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__clkbuf_1
X_10276_ rbzero.tex_b1\[61\] rbzero.tex_b1\[62\] _03199_ vssd1 vssd1 vccd1 vccd1 _03200_
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12015_ _04779_ net65 _04786_ _04787_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__a211o_1
XFILLER_78_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17872_ _02129_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__inv_2
XFILLER_94_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19611_ clknet_leaf_53_i_clk _00542_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16823_ _09354_ _09395_ vssd1 vssd1 vccd1 vccd1 _09430_ sky130_fd_sc_hd__and2_1
XFILLER_93_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19542_ clknet_leaf_11_i_clk _00473_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.wall\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16754_ _09014_ _09016_ _09035_ _09036_ vssd1 vssd1 vccd1 vccd1 _09362_ sky130_fd_sc_hd__or4_1
XFILLER_171_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13966_ _06572_ _06587_ _05349_ vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__mux2_1
XFILLER_185_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15705_ _08386_ _08387_ vssd1 vssd1 vccd1 vccd1 _08388_ sky130_fd_sc_hd__and2_1
X_12917_ _05671_ _05672_ _05673_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__o21a_1
X_16685_ _09130_ _09180_ _09178_ vssd1 vssd1 vccd1 vccd1 _09294_ sky130_fd_sc_hd__a21oi_1
XFILLER_46_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19473_ clknet_leaf_51_i_clk _00419_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13897_ _05325_ _06602_ _06651_ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__a21o_1
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15636_ _07011_ _08317_ _08318_ vssd1 vssd1 vccd1 vccd1 _08319_ sky130_fd_sc_hd__a21o_1
X_12848_ _05586_ _05598_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__nor2_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15567_ _08246_ _08248_ _08250_ vssd1 vssd1 vccd1 vccd1 _08251_ sky130_fd_sc_hd__o21ai_1
X_18355_ rbzero.pov.sclk_buffer\[2\] rbzero.pov.sclk_buffer\[1\] vssd1 vssd1 vccd1
+ vccd1 _02414_ sky130_fd_sc_hd__nor2b_2
X_12779_ _05404_ _05425_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__xnor2_4
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518_ _07189_ _07205_ vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__nor2_1
X_17306_ _01628_ _01629_ _01630_ vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__o21ai_1
XFILLER_148_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15498_ _08174_ _08175_ _08177_ vssd1 vssd1 vccd1 vccd1 _08182_ sky130_fd_sc_hd__a21oi_1
X_18286_ _02375_ vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14449_ _07136_ vssd1 vssd1 vccd1 vccd1 _07137_ sky130_fd_sc_hd__clkbuf_4
X_17237_ rbzero.wall_tracer.trackDistY\[-3\] rbzero.wall_tracer.stepDistY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__nor2_1
XFILLER_190_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17168_ _01458_ _01511_ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__xnor2_4
X_16119_ _08731_ vssd1 vssd1 vccd1 vccd1 _08732_ sky130_fd_sc_hd__inv_2
XFILLER_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17099_ _09629_ _09609_ _09703_ vssd1 vssd1 vccd1 vccd1 _09704_ sky130_fd_sc_hd__a21o_1
X_09990_ rbzero.tex_r0\[5\] rbzero.tex_r0\[4\] _03039_ vssd1 vssd1 vccd1 vccd1 _03049_
+ sky130_fd_sc_hd__mux2_1
XFILLER_192_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19809_ clknet_leaf_15_i_clk _00740_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19208__366 clknet_1_1__leaf__02751_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__inv_2
XFILLER_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20515_ clknet_leaf_79_i_clk _01446_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20446_ net506 _01377_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20377_ net437 _01308_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_192_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10130_ rbzero.tex_g1\[2\] rbzero.tex_g1\[3\] _03117_ vssd1 vssd1 vccd1 vccd1 _03123_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10061_ rbzero.tex_g1\[35\] rbzero.tex_g1\[36\] _03084_ vssd1 vssd1 vccd1 vccd1 _03087_
+ sky130_fd_sc_hd__mux2_1
XFILLER_121_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13820_ _06197_ _06216_ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__and2_1
XFILLER_29_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13751_ _06478_ _06505_ _06507_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__a21bo_1
X_10963_ _03747_ _03748_ _03693_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__mux2_1
XFILLER_189_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12702_ _05270_ _05441_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__or2_1
XFILLER_71_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16470_ _09076_ _09079_ _09080_ vssd1 vssd1 vccd1 vccd1 _09081_ sky130_fd_sc_hd__a21oi_4
X_13682_ _05527_ _06071_ vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__nor2_1
X_10894_ _03674_ _03678_ _03679_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__a21o_1
XFILLER_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15421_ _08104_ _08105_ vssd1 vssd1 vccd1 vccd1 _08106_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12633_ _05369_ _05334_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__nand2_4
XFILLER_31_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15352_ _07874_ _07913_ _08037_ vssd1 vssd1 vccd1 vccd1 _08038_ sky130_fd_sc_hd__a21oi_1
XFILLER_12_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18140_ _02282_ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__buf_2
XFILLER_19_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12564_ _05269_ _05320_ vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14303_ _06989_ _06990_ _06914_ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__mux2_1
X_11515_ rbzero.tex_g1\[43\] rbzero.tex_g1\[42\] _03727_ vssd1 vssd1 vccd1 vccd1 _04298_
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18071_ _02239_ vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__clkbuf_1
X_15283_ _07859_ _07868_ _07867_ vssd1 vssd1 vccd1 vccd1 _07969_ sky130_fd_sc_hd__a21o_1
XFILLER_89_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12495_ _05202_ _05203_ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__nand2_1
XFILLER_89_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17022_ _09626_ _09627_ _08507_ vssd1 vssd1 vccd1 vccd1 _09628_ sky130_fd_sc_hd__o21a_1
XFILLER_156_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14234_ rbzero.debug_overlay.playerY\[-6\] _06877_ vssd1 vssd1 vccd1 vccd1 _06922_
+ sky130_fd_sc_hd__or2_1
XFILLER_156_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11446_ _04150_ _04229_ _03830_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__mux2_1
XFILLER_165_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14165_ _06852_ vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__buf_4
X_11377_ rbzero.tex_g0\[25\] rbzero.tex_g0\[24\] _03709_ vssd1 vssd1 vccd1 vccd1 _04161_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13116_ _05859_ _05860_ _05872_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__a21o_1
X_10328_ rbzero.tex_b1\[36\] rbzero.tex_b1\[37\] _03221_ vssd1 vssd1 vccd1 vccd1 _03227_
+ sky130_fd_sc_hd__mux2_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14096_ rbzero.wall_tracer.trackDistY\[8\] _06785_ _06811_ vssd1 vssd1 vccd1 vccd1
+ _00447_ sky130_fd_sc_hd__o21a_1
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ _02161_ vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__clkbuf_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _05779_ _05803_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__xnor2_1
XFILLER_59_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10259_ rbzero.tex_g0\[6\] rbzero.tex_g0\[5\] _03188_ vssd1 vssd1 vccd1 vccd1 _03191_
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19235__10 clknet_1_1__leaf__02754_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__inv_2
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17855_ rbzero.spi_registers.spi_counter\[2\] _02115_ vssd1 vssd1 vccd1 vccd1 _02116_
+ sky130_fd_sc_hd__nand2_1
XFILLER_120_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16806_ _09410_ _09413_ vssd1 vssd1 vccd1 vccd1 _09414_ sky130_fd_sc_hd__nand2_1
XFILLER_93_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19250__24 clknet_1_1__leaf__02755_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__inv_2
X_17786_ _02050_ _02051_ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__nand2_1
XFILLER_54_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14998_ _07648_ _07667_ _07685_ vssd1 vssd1 vccd1 vccd1 _07686_ sky130_fd_sc_hd__o21a_1
X_19525_ clknet_leaf_49_i_clk _00471_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16737_ _09335_ _09344_ vssd1 vssd1 vccd1 vccd1 _09345_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13949_ _05324_ _06620_ _06639_ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__o21ai_1
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19456_ clknet_leaf_35_i_clk _00402_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16668_ _09268_ _09276_ vssd1 vssd1 vccd1 vccd1 _09277_ sky130_fd_sc_hd__nand2_1
XFILLER_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15619_ _08299_ _08302_ vssd1 vssd1 vccd1 vccd1 _08303_ sky130_fd_sc_hd__xor2_4
X_19387_ _08439_ _02862_ _02863_ _02319_ rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1
+ _01426_ sky130_fd_sc_hd__a32o_1
X_16599_ _09127_ _09205_ _09207_ vssd1 vssd1 vccd1 vccd1 _09208_ sky130_fd_sc_hd__a21oi_1
XFILLER_15_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18338_ _02404_ vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18269_ rbzero.spi_registers.spi_buffer\[4\] rbzero.spi_registers.new_sky\[4\] _02361_
+ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__mux2_1
XFILLER_163_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20300_ net360 _01231_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20231_ net291 _01162_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20162_ net222 _01093_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[9\] sky130_fd_sc_hd__dfxtp_1
X_09973_ _03040_ vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20093_ clknet_leaf_8_i_clk _01024_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18419__60 clknet_1_1__leaf__02437_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__inv_2
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18434__74 clknet_1_0__leaf__02438_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__inv_2
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18924__109 clknet_1_0__leaf__02724_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__inv_2
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11300_ _04058_ _04070_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__nor2_4
XFILLER_126_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12280_ _05035_ _05036_ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__and2_1
XFILLER_5_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11231_ gpout0.vpos\[6\] _03838_ _04008_ _04015_ vssd1 vssd1 vccd1 vccd1 _04016_
+ sky130_fd_sc_hd__or4_1
X_20429_ net489 _01360_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11162_ rbzero.tex_r1\[40\] _03920_ _03618_ _03945_ _03946_ vssd1 vssd1 vccd1 vccd1
+ _03947_ sky130_fd_sc_hd__a311o_1
XFILLER_134_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10113_ rbzero.tex_g1\[10\] rbzero.tex_g1\[11\] _03106_ vssd1 vssd1 vccd1 vccd1 _03114_
+ sky130_fd_sc_hd__mux2_1
X_11093_ _03517_ rbzero.map_overlay.i_othery\[0\] vssd1 vssd1 vccd1 vccd1 _03879_
+ sky130_fd_sc_hd__nand2_1
X_15970_ _08584_ vssd1 vssd1 vccd1 vccd1 _08585_ sky130_fd_sc_hd__inv_2
XFILLER_150_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14921_ _07575_ _07576_ _07608_ vssd1 vssd1 vccd1 vccd1 _07609_ sky130_fd_sc_hd__and3_1
X_10044_ rbzero.tex_g1\[43\] rbzero.tex_g1\[44\] _03073_ vssd1 vssd1 vccd1 vccd1 _03078_
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17640_ _04100_ rbzero.wall_tracer.rayAddendX\[-5\] vssd1 vssd1 vccd1 vccd1 _01917_
+ sky130_fd_sc_hd__nand2_1
XFILLER_76_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14852_ _06865_ _06968_ vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__or2_1
XFILLER_60_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13803_ _06435_ _06470_ _06430_ _06472_ _06559_ vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__a32o_1
X_17571_ _01855_ _01856_ _01853_ _01854_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__o211ai_2
XFILLER_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14783_ _07427_ _07470_ vssd1 vssd1 vccd1 vccd1 _07471_ sky130_fd_sc_hd__nor2_1
X_11995_ net31 _04768_ net32 vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__or3b_1
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19310_ _02794_ _02795_ _02797_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__o21ai_1
X_16522_ _09031_ _09044_ vssd1 vssd1 vccd1 vccd1 _09132_ sky130_fd_sc_hd__nand2_1
X_13734_ _06455_ _06487_ _06488_ _06490_ vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__a22o_1
XFILLER_1_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10946_ _03662_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__buf_4
XFILLER_17_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16453_ _09061_ _09062_ vssd1 vssd1 vccd1 vccd1 _09064_ sky130_fd_sc_hd__nand2_1
X_13665_ _06399_ _06420_ _06421_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__a21o_1
X_10877_ _03662_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__buf_4
XFILLER_143_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _08088_ _07948_ _07951_ vssd1 vssd1 vccd1 vccd1 _08089_ sky130_fd_sc_hd__o21a_1
X_12616_ _05335_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__clkbuf_4
X_16384_ _08993_ _08994_ vssd1 vssd1 vccd1 vccd1 _08995_ sky130_fd_sc_hd__nor2_1
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _06232_ _06352_ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__or2_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15335_ _07898_ _08020_ vssd1 vssd1 vccd1 vccd1 _08021_ sky130_fd_sc_hd__and2_1
XFILLER_118_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18123_ rbzero.spi_registers.new_other\[10\] _02264_ _02271_ _02266_ vssd1 vssd1
+ vccd1 vccd1 _00754_ sky130_fd_sc_hd__o211a_1
XFILLER_185_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12547_ _05303_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__buf_2
XFILLER_185_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15266_ _07950_ _07949_ vssd1 vssd1 vccd1 vccd1 _07952_ sky130_fd_sc_hd__or2b_1
X_18054_ rbzero.spi_registers.spi_buffer\[3\] rbzero.spi_registers.spi_buffer\[2\]
+ _02227_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__mux2_1
X_12478_ _05120_ _05234_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__or2_2
XANTENNA_3 _04150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17005_ _09609_ _09610_ vssd1 vssd1 vccd1 vccd1 _09611_ sky130_fd_sc_hd__nand2_1
X_14217_ _06852_ _06712_ _06904_ _06859_ vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__o211a_2
X_11429_ _03656_ _04210_ _04212_ _03669_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__o211a_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15197_ _07882_ _07883_ vssd1 vssd1 vccd1 vccd1 _07884_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14148_ _03389_ _03454_ vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__and2_1
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14079_ rbzero.wall_tracer.visualWallDist\[0\] _06796_ _06785_ rbzero.wall_tracer.trackDistY\[0\]
+ _06797_ vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__o221a_1
XFILLER_141_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17907_ _02152_ vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__clkbuf_1
X_18887_ _03902_ _04503_ _02280_ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__and3_1
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17838_ _01972_ _02085_ _03340_ _02094_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__o211a_1
XFILLER_39_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17769_ _02036_ vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19508_ clknet_leaf_56_i_clk _00454_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19439_ gpout2.clk_div\[0\] gpout2.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__nand2_1
XFILLER_179_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20214_ net274 _01145_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09956_ _03031_ vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__clkbuf_1
X_20145_ clknet_leaf_12_i_clk _01076_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[3\] sky130_fd_sc_hd__dfxtp_4
XFILLER_104_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09887_ _02983_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__clkbuf_4
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20076_ clknet_leaf_8_i_clk _01007_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10800_ rbzero.traced_texVinit\[6\] rbzero.spi_registers.vshift\[3\] vssd1 vssd1
+ vccd1 vccd1 _03586_ sky130_fd_sc_hd__nand2_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ net19 _04555_ _04556_ net18 vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__a31o_1
XFILLER_198_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10731_ gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__clkbuf_4
XFILLER_201_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13450_ _06079_ _06139_ _06206_ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__a21oi_1
XFILLER_201_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10662_ _03341_ _03457_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__or2_4
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12401_ _05154_ _05157_ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__xnor2_2
XFILLER_90_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13381_ _06118_ _06137_ _06135_ vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__a21oi_1
XFILLER_167_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10593_ _03368_ _03383_ _03387_ _03388_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__o211a_1
XFILLER_166_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15120_ _07703_ _07807_ vssd1 vssd1 vccd1 vccd1 _07808_ sky130_fd_sc_hd__xor2_4
X_12332_ _03479_ _04909_ _04910_ _05088_ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__a31o_1
XFILLER_194_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15051_ _07731_ _07737_ vssd1 vssd1 vccd1 vccd1 _07739_ sky130_fd_sc_hd__or2_1
X_12263_ _05019_ _05020_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__nand2_1
XFILLER_107_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14002_ _05373_ _06740_ _06745_ _05476_ _06629_ vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__a221o_4
X_11214_ _03638_ _03643_ _03998_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__o21a_1
XFILLER_123_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12194_ rbzero.wall_tracer.trackDistY\[8\] vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__inv_2
XFILLER_122_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18810_ _02637_ vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__clkbuf_4
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 o_rgb[14] sky130_fd_sc_hd__buf_2
X_11145_ rbzero.tex_r1\[62\] _03767_ vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__or2_1
XFILLER_123_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19790_ clknet_leaf_7_i_clk _00721_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18741_ rbzero.debug_overlay.playerY\[3\] _02614_ _02412_ vssd1 vssd1 vccd1 vccd1
+ _02621_ sky130_fd_sc_hd__a21o_1
XFILLER_89_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11076_ rbzero.map_overlay.i_mapdx\[2\] _03460_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__xor2_1
X_15953_ rbzero.wall_tracer.trackDistX\[-3\] rbzero.wall_tracer.stepDistX\[-3\] vssd1
+ vssd1 vccd1 vccd1 _08570_ sky130_fd_sc_hd__nor2_1
XFILLER_48_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10027_ _03068_ vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__clkbuf_1
X_14904_ _07590_ _07591_ vssd1 vssd1 vccd1 vccd1 _07592_ sky130_fd_sc_hd__nand2_1
XFILLER_37_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18672_ _02566_ _02567_ _02535_ vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__a21oi_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15884_ rbzero.wall_tracer.state\[1\] vssd1 vssd1 vccd1 vccd1 _08509_ sky130_fd_sc_hd__buf_8
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17623_ _04933_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__inv_2
XFILLER_63_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14835_ _07498_ _07521_ vssd1 vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__nor2_1
XFILLER_63_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18413__55 clknet_1_1__leaf__02436_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__inv_2
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _01785_ rbzero.wall_tracer.rayAddendY\[6\] vssd1 vssd1 vccd1 vccd1 _01842_
+ sky130_fd_sc_hd__xnor2_1
X_11978_ net29 _04751_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__nand2_1
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14766_ _07449_ _07452_ _07453_ vssd1 vssd1 vccd1 vccd1 _07454_ sky130_fd_sc_hd__a21oi_1
X_16505_ _09113_ _09114_ vssd1 vssd1 vccd1 vccd1 _09115_ sky130_fd_sc_hd__and2_1
X_10929_ _03583_ _03582_ _03598_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__nor3_1
X_13717_ _06436_ _06473_ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__and2_1
X_17485_ rbzero.debug_overlay.vplaneY\[-3\] rbzero.debug_overlay.vplaneY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__and2_1
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14697_ _06900_ _07147_ vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__nor2_1
XFILLER_149_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16436_ _07661_ _07662_ vssd1 vssd1 vccd1 vccd1 _09047_ sky130_fd_sc_hd__and2_1
X_13648_ _06385_ _06386_ _06387_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__a21oi_1
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16367_ _08976_ _08977_ vssd1 vssd1 vccd1 vccd1 _08978_ sky130_fd_sc_hd__nand2_1
X_13579_ _06297_ _06300_ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_53_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_185_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18106_ _03517_ gpout0.vpos\[2\] gpout0.vpos\[1\] gpout0.vpos\[0\] vssd1 vssd1 vccd1
+ vccd1 _02259_ sky130_fd_sc_hd__and4_1
X_15318_ _07881_ _07994_ _08003_ vssd1 vssd1 vccd1 vccd1 _08004_ sky130_fd_sc_hd__a21o_1
XFILLER_145_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16298_ _08392_ _08799_ _08800_ _08798_ vssd1 vssd1 vccd1 vccd1 _08910_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18037_ _02220_ vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15249_ _06914_ vssd1 vssd1 vccd1 vccd1 _07936_ sky130_fd_sc_hd__inv_2
XFILLER_67_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_68_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09810_ rbzero.tex_r1\[24\] rbzero.tex_r1\[25\] _02943_ vssd1 vssd1 vccd1 vccd1 _02953_
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19988_ clknet_leaf_87_i_clk _00919_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09741_ rbzero.tex_r1\[57\] rbzero.tex_r1\[58\] _02910_ vssd1 vssd1 vccd1 vccd1 _02917_
+ sky130_fd_sc_hd__mux2_1
XFILLER_140_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__02439_ clknet_0__02439_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02439_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_55_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20128_ clknet_leaf_78_i_clk _01059_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09939_ _03022_ vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12950_ _05704_ _05705_ _05706_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__nand3_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20059_ clknet_leaf_0_i_clk _00990_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.mosi sky130_fd_sc_hd__dfxtp_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901_ _04670_ _04675_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__nand2_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _05520_ _05521_ _05637_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__o21ai_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14620_ _07293_ _07307_ vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__xnor2_1
X_11832_ _04595_ _04601_ _04608_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__or3b_2
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _07223_ _07224_ _07238_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__a21o_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _03464_ _04512_ _04516_ _03474_ _04496_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__a221o_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13502_ _06239_ _06258_ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__xnor2_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ gpout0.hpos\[2\] _03501_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__nand2_1
XFILLER_201_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _06759_ _07165_ vssd1 vssd1 vccd1 vccd1 _07170_ sky130_fd_sc_hd__nand2_1
X_17270_ _01534_ _01599_ _01600_ _01526_ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__a31o_1
X_11694_ _03838_ _03465_ _04019_ _03529_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__nand4_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16221_ _08832_ _08833_ vssd1 vssd1 vccd1 vccd1 _08834_ sky130_fd_sc_hd__xnor2_4
X_13433_ _06188_ _06189_ vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__nor2_1
XFILLER_201_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10645_ rbzero.map_overlay.i_otherx\[4\] vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__inv_2
XFILLER_155_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16152_ _08661_ _08670_ vssd1 vssd1 vccd1 vccd1 _08765_ sky130_fd_sc_hd__or2b_1
XFILLER_139_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13364_ _05551_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__buf_2
XFILLER_6_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10576_ _03370_ _03371_ rbzero.wall_tracer.mapY\[7\] vssd1 vssd1 vccd1 vccd1 _03372_
+ sky130_fd_sc_hd__a21o_1
X_15103_ _07783_ _07789_ vssd1 vssd1 vccd1 vccd1 _07791_ sky130_fd_sc_hd__or2_1
X_12315_ rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__inv_2
XFILLER_181_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16083_ _08660_ _08696_ vssd1 vssd1 vccd1 vccd1 _08697_ sky130_fd_sc_hd__xnor2_2
XFILLER_182_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13295_ _05982_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__inv_2
XFILLER_6_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15034_ _07720_ _07721_ vssd1 vssd1 vccd1 vccd1 _07722_ sky130_fd_sc_hd__nor2_1
X_19911_ clknet_leaf_19_i_clk _00842_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_vinf
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12246_ _04930_ _04944_ _04926_ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__o21ai_1
XFILLER_170_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19842_ clknet_leaf_18_i_clk _00773_ vssd1 vssd1 vccd1 vccd1 rbzero.mapdxw\[0\] sky130_fd_sc_hd__dfxtp_1
X_12177_ _04937_ _04938_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__nor2_1
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11128_ _03913_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__inv_2
X_19773_ clknet_leaf_5_i_clk _00704_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16985_ _09589_ _09590_ vssd1 vssd1 vccd1 vccd1 _09591_ sky130_fd_sc_hd__xor2_1
XFILLER_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18724_ net40 net39 vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__nor2_1
XFILLER_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11059_ rbzero.debug_overlay.playerX\[4\] _02901_ vssd1 vssd1 vccd1 vccd1 _03845_
+ sky130_fd_sc_hd__xor2_1
XFILLER_77_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15936_ rbzero.wall_tracer.trackDistX\[-5\] rbzero.wall_tracer.stepDistX\[-5\] vssd1
+ vssd1 vccd1 vccd1 _08555_ sky130_fd_sc_hd__nor2_1
XFILLER_3_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19048__221 clknet_1_1__leaf__02736_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__inv_2
X_18655_ rbzero.pov.ready_buffer\[66\] _07021_ _02539_ vssd1 vssd1 vccd1 vccd1 _02555_
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15867_ rbzero.wall_tracer.mapX\[7\] rbzero.wall_tracer.mapX\[6\] _07825_ vssd1 vssd1
+ vccd1 vccd1 _08495_ sky130_fd_sc_hd__o21a_1
XFILLER_92_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17606_ _01786_ rbzero.wall_tracer.rayAddendY\[10\] vssd1 vssd1 vccd1 vccd1 _01890_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_64_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14818_ _06899_ _07156_ _07177_ _06939_ vssd1 vssd1 vccd1 vccd1 _07506_ sky130_fd_sc_hd__o22a_1
XFILLER_149_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18586_ _02512_ vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15798_ rbzero.row_render.texu\[1\] _08456_ _08453_ rbzero.wall_tracer.texu\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__a22o_1
XFILLER_17_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17537_ _01826_ vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__clkbuf_1
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14749_ _07394_ _07435_ _07436_ vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__a21oi_1
XFILLER_178_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17468_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.debug_overlay.vplaneY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__or2_1
XFILLER_33_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16419_ _09006_ _09029_ vssd1 vssd1 vccd1 vccd1 _09030_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17399_ rbzero.wall_tracer.mapX\[5\] _01698_ _08506_ vssd1 vssd1 vccd1 vccd1 _01699_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19094__263 clknet_1_0__leaf__02740_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__inv_2
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09724_ net46 net45 vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__xor2_4
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10430_ _03143_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__clkbuf_4
XFILLER_183_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10361_ _03244_ vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12100_ _04859_ _04860_ _04861_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__o21ai_1
XFILLER_152_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13080_ _05767_ _05797_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__nand2_1
X_10292_ rbzero.tex_b1\[53\] rbzero.tex_b1\[54\] _03199_ vssd1 vssd1 vccd1 vccd1 _03208_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12031_ gpout0.hpos\[0\] _03527_ _03526_ _04020_ _04790_ net34 vssd1 vssd1 vccd1
+ vccd1 _04804_ sky130_fd_sc_hd__mux4_1
XFILLER_137_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16770_ _08247_ _08245_ _08803_ vssd1 vssd1 vccd1 vccd1 _09378_ sky130_fd_sc_hd__a21oi_1
X_13982_ _06598_ _06600_ _06588_ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__mux2_1
X_15721_ _07673_ _08144_ _08272_ vssd1 vssd1 vccd1 vccd1 _08404_ sky130_fd_sc_hd__and3_1
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ _05467_ _05483_ _05516_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__a21oi_1
XFILLER_58_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15652_ _08332_ _08334_ vssd1 vssd1 vccd1 vccd1 _08335_ sky130_fd_sc_hd__xnor2_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _05491_ _05499_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__nand2_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _07246_ _07290_ vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__xnor2_2
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371_ rbzero.pov.spi_counter\[4\] rbzero.pov.spi_counter\[3\] _02423_ vssd1 vssd1
+ vccd1 vccd1 _02426_ sky130_fd_sc_hd__and3_1
XFILLER_57_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ net17 _04588_ _04591_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__a21o_1
X_12795_ _05491_ _05549_ _05551_ _05392_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _06771_ _06776_ _08266_ _07893_ vssd1 vssd1 vccd1 vccd1 _08267_ sky130_fd_sc_hd__nand4_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _04956_ _01527_ _01645_ vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__a21oi_1
XFILLER_183_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14534_ _06917_ _07092_ vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__or2_1
X_11746_ _04514_ _04518_ _04523_ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__or3_2
XFILLER_183_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17253_ _01578_ _01580_ _01579_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__a21boi_1
X_11677_ _03607_ _04453_ _04457_ _03624_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__a211o_1
XFILLER_128_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14465_ _06860_ rbzero.wall_tracer.stepDistY\[2\] _04840_ vssd1 vssd1 vccd1 vccd1
+ _07153_ sky130_fd_sc_hd__o21a_1
XFILLER_186_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16204_ _08815_ _08816_ vssd1 vssd1 vccd1 vccd1 _08817_ sky130_fd_sc_hd__nand2_1
X_13416_ _06172_ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__clkbuf_2
X_10628_ rbzero.map_overlay.i_mapdx\[2\] _03353_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__xnor2_1
X_14396_ _06940_ vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__buf_2
X_17184_ _01526_ vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__buf_4
XFILLER_183_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16135_ _08746_ _08747_ vssd1 vssd1 vccd1 vccd1 _08748_ sky130_fd_sc_hd__xnor2_1
X_13347_ _06001_ _06060_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__or2_1
XFILLER_183_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10559_ rbzero.debug_overlay.playerY\[0\] _03352_ _03354_ rbzero.debug_overlay.playerX\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16066_ _07213_ _08678_ vssd1 vssd1 vccd1 vccd1 _08680_ sky130_fd_sc_hd__or2_1
XFILLER_143_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13278_ _06002_ _06034_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__xnor2_4
XFILLER_142_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15017_ _07127_ _07086_ vssd1 vssd1 vccd1 vccd1 _07705_ sky130_fd_sc_hd__or2b_1
X_12229_ _04987_ _04988_ _04989_ _04990_ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__and4b_1
XFILLER_142_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19825_ clknet_leaf_14_i_clk _00756_ vssd1 vssd1 vccd1 vccd1 rbzero.map_overlay.i_othery\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19756_ clknet_leaf_88_i_clk _00687_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16968_ _09570_ _09572_ vssd1 vssd1 vccd1 vccd1 _09574_ sky130_fd_sc_hd__and2_1
XFILLER_110_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18707_ rbzero.debug_overlay.playerY\[-6\] _02588_ _02595_ _02586_ vssd1 vssd1 vccd1
+ vccd1 _01014_ sky130_fd_sc_hd__o211a_1
XFILLER_77_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15919_ rbzero.wall_tracer.trackDistX\[-7\] rbzero.wall_tracer.stepDistX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _08540_ sky130_fd_sc_hd__nor2_1
X_19687_ clknet_leaf_68_i_clk _00618_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16899_ _09429_ _09430_ _09504_ vssd1 vssd1 vccd1 vccd1 _09506_ sky130_fd_sc_hd__or3_1
XFILLER_80_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18638_ rbzero.debug_overlay.playerX\[-8\] _02543_ vssd1 vssd1 vccd1 vccd1 _02544_
+ sky130_fd_sc_hd__or2_1
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18569_ _02503_ vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19102__270 clknet_1_0__leaf__02741_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__inv_2
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20462_ net142 _01393_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18959__141 clknet_1_1__leaf__02727_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__inv_2
XFILLER_146_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20393_ net453 _01324_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11600_ _04375_ _04378_ _04381_ _03607_ _03627_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__a221o_1
XFILLER_30_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12580_ _05244_ _05276_ _05297_ _05192_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__a31o_1
XFILLER_70_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11531_ _03522_ _04313_ _04148_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__o21ai_4
XFILLER_157_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14250_ _04838_ rbzero.wall_tracer.stepDistX\[-5\] _06934_ _06937_ vssd1 vssd1 vccd1
+ vccd1 _06938_ sky130_fd_sc_hd__o22ai_4
X_11462_ _04243_ _04244_ _03740_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__mux2_1
XFILLER_165_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13201_ _05952_ _05956_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__and2_1
XFILLER_165_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10413_ _03271_ vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14181_ _04831_ _06868_ _06859_ vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__o21a_1
X_11393_ rbzero.tex_g0\[13\] rbzero.tex_g0\[12\] _03662_ vssd1 vssd1 vccd1 vccd1 _04177_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13132_ _05628_ _05858_ _05887_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__nand3_1
X_10344_ _03235_ vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13063_ _05488_ _05810_ _05812_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__a21bo_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17940_ rbzero.pov.spi_buffer\[24\] rbzero.pov.ready_buffer\[24\] _02164_ vssd1 vssd1
+ vccd1 vccd1 _02170_ sky130_fd_sc_hd__mux2_1
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10275_ _03072_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__clkbuf_4
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12014_ net36 net37 vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__nand2_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17871_ rbzero.spi_registers.spi_counter\[3\] rbzero.spi_registers.spi_counter\[2\]
+ _02112_ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__and3_1
XFILLER_78_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19610_ clknet_leaf_53_i_clk _00541_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
X_16822_ _09393_ _09394_ vssd1 vssd1 vccd1 vccd1 _09429_ sky130_fd_sc_hd__nor2_1
XFILLER_120_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19541_ clknet_leaf_19_i_clk _00472_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.wall\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16753_ _09359_ _09360_ vssd1 vssd1 vccd1 vccd1 _09361_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13965_ _06713_ vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15704_ _08250_ _08378_ _08385_ vssd1 vssd1 vccd1 vccd1 _08387_ sky130_fd_sc_hd__nand3_1
XFILLER_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12916_ _05670_ _05666_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__or2b_1
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19472_ clknet_leaf_51_i_clk _00418_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16684_ _09245_ _09292_ vssd1 vssd1 vccd1 vccd1 _09293_ sky130_fd_sc_hd__xnor2_1
X_13896_ _05367_ _06605_ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__and2_1
X_15635_ _08199_ _08314_ vssd1 vssd1 vccd1 vccd1 _08318_ sky130_fd_sc_hd__xor2_1
XFILLER_61_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12847_ _05583_ _05585_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__and2_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ rbzero.pov.spi_done rbzero.pov.ready _02285_ _02413_ vssd1 vssd1 vccd1 vccd1
+ _00843_ sky130_fd_sc_hd__o211a_1
X_15566_ _07581_ _07198_ _08249_ vssd1 vssd1 vccd1 vccd1 _08250_ sky130_fd_sc_hd__or3_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383__27 clknet_1_0__leaf__02434_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__inv_2
XFILLER_15_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12778_ _05534_ _05515_ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__xnor2_2
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _01628_ _01629_ _01630_ vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__or3_1
X_14517_ _07191_ _07203_ _07204_ vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__a21oi_1
X_11729_ gpout0.vpos\[2\] vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__clkbuf_4
X_18285_ rbzero.spi_registers.spi_buffer\[4\] rbzero.spi_registers.new_floor\[4\]
+ _02370_ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__mux2_1
XFILLER_175_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15497_ rbzero.wall_tracer.texu\[3\] _06853_ _08180_ _08181_ _03498_ vssd1 vssd1
+ vccd1 vccd1 _00478_ sky130_fd_sc_hd__o221a_1
XFILLER_175_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17236_ rbzero.wall_tracer.trackDistY\[-4\] _01558_ _01571_ _08561_ vssd1 vssd1 vccd1
+ vccd1 _00567_ sky130_fd_sc_hd__o22a_1
XFILLER_80_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14448_ _04949_ rbzero.wall_tracer.stepDistX\[1\] _07134_ _07135_ vssd1 vssd1 vccd1
+ vccd1 _07136_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17167_ _01460_ _01510_ vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__xnor2_4
XFILLER_122_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14379_ _06871_ _07037_ _07048_ _07024_ vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__o22a_1
XFILLER_115_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16118_ _07235_ _07972_ _07959_ _08069_ vssd1 vssd1 vccd1 vccd1 _08731_ sky130_fd_sc_hd__or4_1
XFILLER_143_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17098_ _09529_ _09702_ vssd1 vssd1 vccd1 vccd1 _09703_ sky130_fd_sc_hd__xnor2_1
XFILLER_182_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16049_ _07581_ _07530_ _07756_ _07757_ vssd1 vssd1 vccd1 vccd1 _08663_ sky130_fd_sc_hd__or4_1
XFILLER_143_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19808_ clknet_leaf_3_i_clk _00739_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19739_ clknet_leaf_76_i_clk _00670_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20514_ clknet_leaf_77_i_clk _01445_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20445_ net505 _01376_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20376_ net436 _01307_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10060_ _03086_ vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10962_ rbzero.tex_r0\[59\] rbzero.tex_r0\[58\] _03690_ vssd1 vssd1 vccd1 vccd1 _03748_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13750_ _06500_ _06506_ vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__or2b_1
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12701_ _05454_ _05455_ _05457_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__nor3b_2
XFILLER_44_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10893_ _03624_ vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__buf_6
X_13681_ _06399_ _06437_ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15420_ _07735_ _07281_ vssd1 vssd1 vccd1 vccd1 _08105_ sky130_fd_sc_hd__or2_1
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12632_ _05376_ _05388_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__nor2_1
XFILLER_19_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15351_ _07910_ _07912_ vssd1 vssd1 vccd1 vccd1 _08037_ sky130_fd_sc_hd__nor2_1
X_12563_ _05319_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__clkbuf_4
XFILLER_197_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11514_ _04198_ _04292_ _04296_ _03648_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__a211o_1
X_14302_ rbzero.debug_overlay.playerX\[-3\] vssd1 vssd1 vccd1 vccd1 _06990_ sky130_fd_sc_hd__inv_2
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18070_ rbzero.spi_registers.spi_buffer\[11\] rbzero.spi_registers.spi_buffer\[10\]
+ _02226_ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__mux2_1
X_15282_ _07966_ _07967_ vssd1 vssd1 vccd1 vccd1 _07968_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12494_ _05224_ _05226_ _05228_ _05247_ _05250_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__o41a_1
XFILLER_184_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17021_ _09623_ _09624_ _09625_ _04946_ vssd1 vssd1 vccd1 vccd1 _09627_ sky130_fd_sc_hd__a31o_1
X_11445_ _03764_ _04186_ _04224_ _04228_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__a31o_1
X_14233_ _06901_ _06918_ _06920_ vssd1 vssd1 vccd1 vccd1 _06921_ sky130_fd_sc_hd__o21ai_2
XFILLER_109_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14164_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__clkbuf_4
X_11376_ _03671_ _04153_ _04159_ _03704_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__a211o_1
XFILLER_153_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10327_ _03226_ vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__clkbuf_1
X_13115_ _05870_ _05871_ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__nand2_1
XFILLER_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14095_ rbzero.wall_tracer.visualWallDist\[8\] _03495_ _05005_ rbzero.wall_tracer.trackDistX\[8\]
+ _03497_ vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__o221a_1
XFILLER_180_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ rbzero.pov.spi_buffer\[16\] rbzero.pov.ready_buffer\[16\] _02153_ vssd1 vssd1
+ vccd1 vccd1 _02161_ sky130_fd_sc_hd__mux2_1
X_13046_ _05781_ _05780_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__or2b_1
X_10258_ _03190_ vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_191_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17854_ rbzero.spi_registers.spi_counter\[3\] _02111_ _02112_ _02114_ vssd1 vssd1
+ vccd1 vccd1 _02115_ sky130_fd_sc_hd__a31o_1
X_10189_ rbzero.tex_g0\[39\] rbzero.tex_g0\[38\] _03144_ vssd1 vssd1 vccd1 vccd1 _03154_
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16805_ _09092_ _09411_ _09412_ vssd1 vssd1 vccd1 vccd1 _09413_ sky130_fd_sc_hd__a21oi_1
X_17785_ _02001_ rbzero.wall_tracer.rayAddendX\[5\] _02040_ vssd1 vssd1 vccd1 vccd1
+ _02051_ sky130_fd_sc_hd__a21o_1
XFILLER_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14997_ _07648_ _07667_ _07684_ vssd1 vssd1 vccd1 vccd1 _07685_ sky130_fd_sc_hd__a21o_1
XFILLER_47_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19524_ clknet_leaf_49_i_clk _00470_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[9\]
+ sky130_fd_sc_hd__dfxtp_2
X_16736_ _09342_ _09343_ vssd1 vssd1 vccd1 vccd1 _09344_ sky130_fd_sc_hd__nor2_1
XFILLER_34_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13948_ _06603_ _06633_ _06660_ _05347_ vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__a211o_1
XFILLER_93_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19455_ clknet_leaf_64_i_clk _00401_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16667_ _09269_ _09275_ vssd1 vssd1 vccd1 vccd1 _09276_ sky130_fd_sc_hd__xor2_1
X_13879_ _06601_ _06598_ _06634_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__a21o_1
XFILLER_201_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15618_ _08051_ _08300_ _08301_ _08172_ vssd1 vssd1 vccd1 vccd1 _08302_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_195_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19386_ _02854_ _02859_ _02860_ _02861_ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__nand4_1
X_16598_ _09105_ _09106_ _09206_ vssd1 vssd1 vccd1 vccd1 _09207_ sky130_fd_sc_hd__o21a_1
XFILLER_50_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18337_ rbzero.spi_registers.new_vshift\[2\] rbzero.spi_registers.spi_buffer\[2\]
+ _02401_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__mux2_1
XFILLER_175_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15549_ _07281_ _07123_ vssd1 vssd1 vccd1 vccd1 _08233_ sky130_fd_sc_hd__or2_1
XFILLER_175_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18268_ _02365_ vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17219_ _01553_ _01554_ _01555_ _04946_ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__a31o_1
XFILLER_128_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18199_ _03337_ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__buf_6
X_20230_ net290 _01161_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20161_ net221 _01092_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[8\] sky130_fd_sc_hd__dfxtp_1
X_09972_ rbzero.tex_r0\[14\] rbzero.tex_r0\[13\] _03039_ vssd1 vssd1 vccd1 vccd1 _03040_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__02739_ clknet_0__02739_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__02739_
+ sky130_fd_sc_hd__clkbuf_16
X_19214__371 clknet_1_1__leaf__02752_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__inv_2
XFILLER_131_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20092_ clknet_leaf_8_i_clk _01023_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11230_ _03834_ _03524_ _03782_ _03849_ _04014_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__a221o_1
XFILLER_101_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20428_ net488 _01359_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11161_ rbzero.tex_r1\[41\] _03919_ _03926_ _03669_ vssd1 vssd1 vccd1 vccd1 _03946_
+ sky130_fd_sc_hd__a31o_1
XFILLER_134_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20359_ net419 _01290_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10112_ _03113_ vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11092_ gpout0.vpos\[7\] _03871_ _03430_ _03524_ _03877_ vssd1 vssd1 vccd1 vccd1
+ _03878_ sky130_fd_sc_hd__a221o_1
XFILLER_1_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14920_ _07583_ _07607_ _07605_ vssd1 vssd1 vccd1 vccd1 _07608_ sky130_fd_sc_hd__a21bo_1
X_10043_ _03077_ vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14851_ _07536_ _07538_ vssd1 vssd1 vccd1 vccd1 _07539_ sky130_fd_sc_hd__xnor2_1
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13802_ _06435_ _06558_ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__and2_1
XFILLER_91_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17570_ _01853_ _01854_ _01855_ _01856_ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__a211o_1
XFILLER_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14782_ _07443_ _07468_ _07469_ vssd1 vssd1 vccd1 vccd1 _07470_ sky130_fd_sc_hd__a21oi_2
X_11994_ _04743_ _04761_ _04767_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16521_ _09013_ _09025_ _09023_ vssd1 vssd1 vccd1 vccd1 _09131_ sky130_fd_sc_hd__a21o_1
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13733_ _06453_ _06489_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__xnor2_1
XFILLER_72_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10945_ rbzero.tex_r0\[43\] _03729_ _03730_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__and3_1
XFILLER_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16452_ _09061_ _09062_ vssd1 vssd1 vccd1 vccd1 _09063_ sky130_fd_sc_hd__nor2_1
X_19042__216 clknet_1_0__leaf__02735_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__inv_2
XFILLER_32_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13664_ _06400_ _06401_ _06419_ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__and3_1
X_10876_ _03614_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__buf_6
X_15403_ _07943_ vssd1 vssd1 vccd1 vccd1 _08088_ sky130_fd_sc_hd__inv_2
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ _05269_ _05338_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__nand2_2
X_16383_ _08992_ _08991_ vssd1 vssd1 vccd1 vccd1 _08994_ sky130_fd_sc_hd__and2b_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13595_ _05990_ _06230_ _06156_ _05472_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__o22a_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18122_ _03441_ _02263_ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__nand2_1
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15334_ _07175_ _04950_ _03493_ _08015_ vssd1 vssd1 vccd1 vccd1 _08020_ sky130_fd_sc_hd__or4_1
XFILLER_61_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12546_ _05301_ _05302_ _05284_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__or3b_1
XFILLER_172_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18053_ _02230_ vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__clkbuf_1
XFILLER_117_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15265_ _07949_ _07950_ vssd1 vssd1 vccd1 vccd1 _07951_ sky130_fd_sc_hd__or2b_1
XFILLER_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12477_ _05233_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__buf_2
XFILLER_32_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17004_ _09426_ _09608_ vssd1 vssd1 vccd1 vccd1 _09610_ sky130_fd_sc_hd__or2_1
XFILLER_144_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ rbzero.wall_tracer.state\[3\] _06903_ vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__nand2_1
X_11428_ _03610_ _04211_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__or2_1
XFILLER_126_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15196_ _06997_ _07123_ vssd1 vssd1 vccd1 vccd1 _07883_ sky130_fd_sc_hd__nor2_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11359_ _03904_ _04134_ _04143_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__and3b_1
XFILLER_113_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14147_ _06838_ vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14078_ rbzero.wall_tracer.trackDistY\[-1\] _06786_ _06802_ vssd1 vssd1 vccd1 vccd1
+ _00438_ sky130_fd_sc_hd__o21a_1
XFILLER_112_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17906_ rbzero.pov.spi_buffer\[8\] rbzero.pov.ready_buffer\[8\] _02143_ vssd1 vssd1
+ vccd1 vccd1 _02152_ sky130_fd_sc_hd__mux2_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13029_ _05777_ _05778_ _05782_ _05783_ _05785_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__a32o_1
XFILLER_140_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18886_ _04503_ _02280_ _02281_ _02285_ vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__o211a_1
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17837_ _02097_ _02098_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17768_ rbzero.wall_tracer.rayAddendX\[4\] _02035_ _03509_ vssd1 vssd1 vccd1 vccd1
+ _02036_ sky130_fd_sc_hd__mux2_1
XFILLER_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16719_ _09215_ _09325_ _09326_ vssd1 vssd1 vccd1 vccd1 _09327_ sky130_fd_sc_hd__o21a_1
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19507_ clknet_leaf_55_i_clk _00453_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17699_ _01961_ _01964_ _01962_ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__a21bo_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19438_ gpout2.clk_div\[0\] net61 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__nor2_1
XFILLER_23_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19369_ rbzero.texV\[6\] _02762_ _02709_ _02848_ vssd1 vssd1 vccd1 vccd1 _01423_
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20213_ net273 _01144_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20144_ clknet_leaf_13_i_clk _01075_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[2\] sky130_fd_sc_hd__dfxtp_1
X_09955_ rbzero.tex_r0\[22\] rbzero.tex_r0\[21\] _03028_ vssd1 vssd1 vccd1 vccd1 _03031_
+ sky130_fd_sc_hd__mux2_1
XFILLER_132_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20075_ clknet_leaf_86_i_clk _01006_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_58_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09886_ _02994_ vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__clkbuf_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10730_ gpout0.vpos\[9\] gpout0.vpos\[8\] _03515_ net2 vssd1 vssd1 vccd1 vccd1 _03516_
+ sky130_fd_sc_hd__or4b_1
XFILLER_41_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10661_ _03389_ _03456_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__nand2_2
XFILLER_90_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12400_ _05155_ _05156_ _05080_ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__o21a_1
XFILLER_167_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13380_ _06135_ _06136_ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__nor2_1
X_10592_ rbzero.wall_tracer.visualWallDist\[10\] vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__inv_2
XFILLER_127_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12331_ rbzero.wall_tracer.visualWallDist\[-2\] _05067_ _03487_ vssd1 vssd1 vccd1
+ vccd1 _05088_ sky130_fd_sc_hd__a21o_1
XFILLER_181_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15050_ _07731_ _07737_ vssd1 vssd1 vccd1 vccd1 _07738_ sky130_fd_sc_hd__nand2_1
XFILLER_5_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12262_ _05019_ _05020_ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__or2_1
XFILLER_108_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11213_ rbzero.row_render.wall\[1\] _03997_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__nand2_1
X_14001_ _06743_ _06744_ _06675_ vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__mux2_1
XFILLER_108_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12193_ _04954_ rbzero.wall_tracer.trackDistX\[9\] vssd1 vssd1 vccd1 vccd1 _04955_
+ sky130_fd_sc_hd__nand2_1
XFILLER_135_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11144_ _03918_ _03922_ _03924_ _03928_ _03721_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__o221a_1
XFILLER_122_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 o_rgb[15] sky130_fd_sc_hd__buf_2
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18740_ _02619_ vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__inv_2
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11075_ rbzero.map_overlay.i_mapdx\[3\] _03838_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__xor2_1
X_15952_ rbzero.wall_tracer.trackDistX\[-3\] vssd1 vssd1 vccd1 vccd1 _08569_ sky130_fd_sc_hd__inv_2
XFILLER_49_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10026_ rbzero.tex_g1\[51\] rbzero.tex_g1\[52\] _03061_ vssd1 vssd1 vccd1 vccd1 _03068_
+ sky130_fd_sc_hd__mux2_1
X_14903_ _06969_ _07157_ _07178_ _06978_ vssd1 vssd1 vccd1 vccd1 _07591_ sky130_fd_sc_hd__o22ai_1
X_18671_ rbzero.debug_overlay.playerX\[1\] _02561_ rbzero.debug_overlay.playerX\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__o21ai_1
XFILLER_48_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15883_ _08507_ vssd1 vssd1 vccd1 vccd1 _08508_ sky130_fd_sc_hd__clkbuf_4
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17622_ _01902_ vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14834_ _07498_ _07521_ vssd1 vssd1 vccd1 vccd1 _07522_ sky130_fd_sc_hd__xor2_1
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17553_ _01745_ _01832_ _01833_ _01841_ vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__a31o_1
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ _07078_ _07178_ _07450_ vssd1 vssd1 vccd1 vccd1 _07453_ sky130_fd_sc_hd__nor3_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11977_ _03906_ _04499_ _03909_ _04500_ _04737_ _04750_ vssd1 vssd1 vccd1 vccd1 _04751_
+ sky130_fd_sc_hd__mux4_1
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16504_ _07878_ _07333_ _07784_ _08767_ vssd1 vssd1 vccd1 vccd1 _09114_ sky130_fd_sc_hd__a2bb2o_1
X_13716_ _06438_ _06468_ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__nand2_1
X_10928_ _03674_ _03708_ _03713_ _03679_ vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__a211o_1
X_17484_ rbzero.debug_overlay.vplaneY\[-3\] rbzero.debug_overlay.vplaneY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__nor2_1
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14696_ _06787_ _04839_ _06985_ _06905_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__and4_1
XFILLER_108_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16435_ _08678_ vssd1 vssd1 vccd1 vccd1 _09046_ sky130_fd_sc_hd__buf_2
XFILLER_20_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13647_ _06373_ _06372_ _06363_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__a21o_1
XFILLER_176_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10859_ _03638_ _03643_ _03644_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__o21a_1
XFILLER_20_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19154_ clknet_1_1__leaf__02743_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__buf_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _08107_ _07960_ _08071_ _07984_ vssd1 vssd1 vccd1 vccd1 _08977_ sky130_fd_sc_hd__o22ai_1
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _06330_ _06334_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__nor2_1
XFILLER_118_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18105_ _03909_ _02257_ _03907_ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__nor3_2
X_15317_ _07995_ _08002_ vssd1 vssd1 vccd1 vccd1 _08003_ sky130_fd_sc_hd__xor2_1
XFILLER_184_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12529_ _05185_ _05208_ _05258_ _05231_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__and4_1
X_16297_ _08791_ _08792_ _08789_ vssd1 vssd1 vccd1 vccd1 _08909_ sky130_fd_sc_hd__a21o_1
XFILLER_145_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18036_ rbzero.pov.spi_buffer\[70\] rbzero.pov.ready_buffer\[70\] _02142_ vssd1 vssd1
+ vccd1 vccd1 _02220_ sky130_fd_sc_hd__mux2_1
X_15248_ _07810_ _07822_ _07933_ vssd1 vssd1 vccd1 vccd1 _07935_ sky130_fd_sc_hd__nand3_1
XFILLER_172_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15179_ _07865_ _07281_ _07716_ _07714_ vssd1 vssd1 vccd1 vccd1 _07866_ sky130_fd_sc_hd__o31a_1
XFILLER_193_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18953__136 clknet_1_0__leaf__02726_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__inv_2
XFILLER_113_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19987_ clknet_leaf_0_i_clk _00918_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09740_ _02916_ vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
.ends

